magic
tech sky130l
timestamp 1753821931
<< nwell >>
rect 5 49 29 62
rect 5 33 39 49
rect 75 45 92 62
rect 75 33 117 45
<< ndiffusion >>
rect 15 27 20 28
rect 15 24 16 27
rect 19 24 20 27
rect 15 22 20 24
rect 22 26 27 28
rect 22 23 23 26
rect 26 23 27 26
rect 22 22 27 23
rect 31 27 36 28
rect 31 24 32 27
rect 35 24 36 27
rect 31 22 36 24
rect 42 27 47 28
rect 42 24 43 27
rect 46 24 47 27
rect 42 22 47 24
rect 69 26 76 28
rect 69 23 71 26
rect 74 23 76 26
rect 69 22 76 23
rect 72 18 76 22
rect 78 18 83 28
rect 85 27 90 28
rect 85 24 86 27
rect 89 24 90 27
rect 85 22 90 24
rect 92 27 97 28
rect 92 24 93 27
rect 96 24 97 27
rect 92 22 97 24
rect 85 18 89 22
<< ndc >>
rect 16 24 19 27
rect 23 23 26 26
rect 32 24 35 27
rect 43 24 46 27
rect 71 23 74 26
rect 86 24 89 27
rect 93 24 96 27
<< ntransistor >>
rect 20 22 22 28
rect 27 22 31 28
rect 47 22 69 28
rect 76 18 78 28
rect 83 18 85 28
rect 90 22 92 28
<< pdiffusion >>
rect 8 56 13 59
rect 8 53 9 56
rect 12 53 13 56
rect 8 36 13 53
rect 15 36 20 59
rect 22 46 26 59
rect 78 56 83 59
rect 78 53 79 56
rect 82 53 83 56
rect 22 41 27 46
rect 22 38 23 41
rect 26 38 27 41
rect 22 36 27 38
rect 31 40 36 46
rect 31 37 32 40
rect 35 37 36 40
rect 31 36 36 37
rect 78 36 83 53
rect 85 42 89 59
rect 85 40 90 42
rect 85 37 86 40
rect 89 37 90 40
rect 85 36 90 37
rect 92 36 95 42
rect 109 41 114 42
rect 109 38 110 41
rect 113 38 114 41
rect 109 36 114 38
<< pdc >>
rect 9 53 12 56
rect 79 53 82 56
rect 23 38 26 41
rect 32 37 35 40
rect 86 37 89 40
rect 110 38 113 41
<< ptransistor >>
rect 13 36 15 59
rect 20 36 22 59
rect 27 36 31 46
rect 83 36 85 59
rect 90 36 92 42
rect 95 36 109 42
<< polysilicon >>
rect 8 66 15 68
rect 8 63 10 66
rect 13 63 15 66
rect 8 61 15 63
rect 13 59 15 61
rect 20 66 27 68
rect 20 63 22 66
rect 25 63 27 66
rect 20 61 27 63
rect 80 66 87 68
rect 80 63 82 66
rect 85 63 87 66
rect 80 61 87 63
rect 20 59 22 61
rect 83 59 85 61
rect 27 53 35 55
rect 27 50 30 53
rect 33 50 35 53
rect 27 48 35 50
rect 27 46 31 48
rect 54 37 61 39
rect 13 34 15 36
rect 20 28 22 36
rect 27 28 31 36
rect 54 34 56 37
rect 59 34 61 37
rect 90 52 99 54
rect 90 49 94 52
rect 97 49 99 52
rect 90 47 99 49
rect 90 42 92 47
rect 95 42 109 44
rect 54 30 61 34
rect 47 28 69 30
rect 76 28 78 30
rect 83 28 85 36
rect 90 28 92 36
rect 95 34 109 36
rect 99 32 106 34
rect 99 29 101 32
rect 104 29 106 32
rect 20 20 22 22
rect 27 20 31 22
rect 47 20 69 22
rect 99 27 106 29
rect 90 20 92 22
rect 76 14 78 18
rect 83 16 85 18
rect 76 12 79 14
rect 77 10 84 12
rect 77 7 79 10
rect 82 7 84 10
rect 77 5 84 7
<< pc >>
rect 10 63 13 66
rect 22 63 25 66
rect 82 63 85 66
rect 30 50 33 53
rect 56 34 59 37
rect 94 49 97 52
rect 101 29 104 32
rect 79 7 82 10
<< m1 >>
rect 8 66 15 68
rect 8 63 10 66
rect 13 63 15 66
rect 8 61 15 63
rect 20 66 27 68
rect 20 63 22 66
rect 25 63 27 66
rect 20 61 27 63
rect 80 66 87 68
rect 80 63 82 66
rect 85 63 87 66
rect 80 61 87 63
rect 9 56 12 58
rect 79 56 82 58
rect 9 51 12 53
rect 28 53 35 55
rect 28 50 30 53
rect 33 50 35 53
rect 79 51 82 53
rect 92 52 99 54
rect 28 48 35 50
rect 92 49 94 52
rect 97 49 99 52
rect 16 27 19 47
rect 92 47 99 49
rect 23 41 26 43
rect 23 36 26 38
rect 32 40 35 42
rect 86 40 89 46
rect 16 22 19 24
rect 23 26 26 28
rect 23 20 26 23
rect 32 27 35 37
rect 54 37 61 39
rect 54 34 56 37
rect 59 34 61 37
rect 54 32 61 34
rect 32 22 35 24
rect 43 27 46 29
rect 43 22 46 24
rect 71 26 74 28
rect 71 17 74 23
rect 86 27 89 37
rect 110 41 113 43
rect 110 36 113 38
rect 99 32 106 34
rect 99 29 101 32
rect 104 29 106 32
rect 86 22 89 24
rect 93 27 96 29
rect 99 27 106 29
rect 93 22 96 24
rect 77 10 84 12
rect 77 7 79 10
rect 82 7 84 10
rect 77 5 84 7
<< m2c >>
rect 10 63 13 66
rect 22 63 25 66
rect 82 63 85 66
rect 9 53 12 56
rect 30 50 33 53
rect 79 53 82 56
rect 16 47 19 50
rect 94 49 97 52
rect 86 46 89 49
rect 23 38 26 41
rect 32 42 35 45
rect 56 34 59 37
rect 43 24 46 27
rect 23 17 26 20
rect 110 38 113 41
rect 101 29 104 32
rect 93 24 96 27
rect 71 14 74 17
rect 79 7 82 10
<< m2 >>
rect 9 66 14 67
rect 9 63 10 66
rect 13 63 14 66
rect 9 62 14 63
rect 21 66 26 67
rect 21 63 22 66
rect 25 63 26 66
rect 21 62 26 63
rect 81 66 86 67
rect 81 63 82 66
rect 85 63 86 66
rect 81 62 86 63
rect 8 56 83 58
rect 8 53 9 56
rect 12 53 13 56
rect 8 52 13 53
rect 29 53 34 54
rect 29 51 30 53
rect 15 50 30 51
rect 33 50 34 53
rect 78 53 79 56
rect 82 53 83 56
rect 78 52 83 53
rect 93 52 98 53
rect 15 47 16 50
rect 19 49 90 50
rect 19 47 20 49
rect 29 48 86 49
rect 15 46 20 47
rect 85 46 86 48
rect 89 46 90 49
rect 31 45 36 46
rect 85 45 90 46
rect 93 49 94 52
rect 97 49 98 52
rect 93 48 98 49
rect 31 42 32 45
rect 35 43 36 45
rect 93 43 95 48
rect 35 42 95 43
rect 22 41 27 42
rect 31 41 95 42
rect 109 41 114 42
rect 22 38 23 41
rect 26 39 27 41
rect 109 39 110 41
rect 26 38 110 39
rect 113 38 114 41
rect 22 37 114 38
rect 55 34 56 37
rect 59 34 60 37
rect 55 33 60 34
rect 100 32 105 33
rect 100 29 101 32
rect 104 29 105 32
rect 100 28 105 29
rect 42 27 47 28
rect 42 24 43 27
rect 46 26 47 27
rect 92 27 97 28
rect 92 26 93 27
rect 46 24 93 26
rect 96 24 97 27
rect 42 23 47 24
rect 92 23 97 24
rect 22 20 27 21
rect 22 17 23 20
rect 26 18 27 20
rect 100 18 102 28
rect 26 17 102 18
rect 22 16 71 17
rect 70 14 71 16
rect 74 16 102 17
rect 74 14 75 16
rect 70 13 75 14
rect 78 10 83 11
rect 78 7 79 10
rect 82 7 83 10
rect 78 6 83 7
<< labels >>
flabel polysilicon 83 31 83 31 3 FreeSerif 8 0 0 0 in(2)
flabel polysilicon 90 31 90 31 3 FreeSerif 8 0 0 0 #10
flabel polysilicon 48 29 48 29 3 FreeSerif 8 0 0 0 Vdd
rlabel polysilicon 13 34 13 34 3 in(1)
rlabel polysilicon 95 34 95 34 3 GND
flabel polysilicon 20 34 20 34 3 FreeSerif 8 0 0 0 in(0)
flabel polysilicon 27 33 27 33 3 FreeSerif 8 0 0 0 out
flabel pdiffusion 8 37 8 37 3 FreeSerif 8 0 0 0 #7
flabel pdiffusion 23 37 23 37 3 FreeSerif 8 0 0 0 Vdd
flabel pdiffusion 32 37 32 37 3 FreeSerif 8 0 0 0 #10
flabel pdiffusion 79 37 79 37 3 FreeSerif 8 0 0 0 #7
flabel pdiffusion 86 37 86 37 3 FreeSerif 8 0 0 0 out
flabel pdiffusion 110 37 110 37 3 FreeSerif 8 0 0 0 Vdd
flabel polysilicon 96 34 96 34 1 FreeSerif 8 0 0 0 GND
flabel ndiffusion 93 23 93 23 3 FreeSerif 8 0 0 0 #12
flabel ndiffusion 86 19 86 19 3 FreeSerif 8 0 0 0 out
flabel polysilicon 76 29 76 29 3 FreeSerif 8 0 0 0 in(3)
flabel ndiffusion 70 23 70 23 3 FreeSerif 8 0 0 0 GND
flabel ndiffusion 43 23 43 23 3 FreeSerif 8 0 0 0 #12
flabel ndiffusion 32 23 32 23 3 FreeSerif 8 0 0 0 #10
flabel ndiffusion 16 23 16 23 3 FreeSerif 8 0 0 0 out
flabel polysilicon 13 35 13 35 3 FreeSerif 8 0 0 0 in(1)
flabel ndiffusion 23 24 23 24 3 FreeSerif 8 0 0 0 GND
flabel m2 11 67 11 67 1 FreeSerif 8 0 0 0 in(1)
port 5 n
flabel m2 24 67 24 67 1 FreeSerif 8 0 0 0 in(0)
port 7 n
flabel m2 83 67 83 67 1 FreeSerif 8 0 0 0 in(2)
port 4 n
flabel m2 s 104 29 105 32 3 FreeSerif 8 0 0 0 GND
port 1 nsew ground input
flabel m2 s 89 46 90 49 3 FreeSerif 8 0 0 0 out
port 6 nsew signal output
flabel m2 s 109 39 110 41 1 FreeSerif 8 0 0 0 Vdd
port 2 nsew power input
flabel m2 83 8 83 8 3 FreeSerif 8 0 0 0 in(3)
port 3 e
rlabel m2 s 25 63 26 66 5 in_50_6
port 1 nsew signal input
rlabel m2 s 22 63 25 66 5 in_50_6
port 1 nsew signal input
rlabel m2 s 21 63 22 66 5 in_50_6
port 1 nsew signal input
rlabel m2 s 21 62 26 63 1 in_50_6
port 1 nsew signal input
rlabel m2 s 21 66 26 67 5 in_50_6
port 1 nsew signal input
rlabel m1 s 25 63 27 66 5 in_50_6
port 1 nsew signal input
rlabel m1 s 22 63 25 66 5 in_50_6
port 1 nsew signal input
rlabel m1 s 20 61 27 63 1 in_50_6
port 1 nsew signal input
rlabel m1 s 20 63 22 66 5 in_50_6
port 1 nsew signal input
rlabel m1 s 20 66 27 68 5 in_50_6
port 1 nsew signal input
rlabel m2 s 13 63 14 66 5 in_51_6
port 2 nsew signal input
rlabel m2 s 10 63 13 66 5 in_51_6
port 2 nsew signal input
rlabel m2 s 9 62 14 63 1 in_51_6
port 2 nsew signal input
rlabel m2 s 9 63 10 66 4 in_51_6
port 2 nsew signal input
rlabel m2 s 9 66 14 67 5 in_51_6
port 2 nsew signal input
rlabel m1 s 13 63 15 66 5 in_51_6
port 2 nsew signal input
rlabel m1 s 10 63 13 66 5 in_51_6
port 2 nsew signal input
rlabel m1 s 8 61 15 63 1 in_51_6
port 2 nsew signal input
rlabel m1 s 8 63 10 66 4 in_51_6
port 2 nsew signal input
rlabel m1 s 8 66 15 68 5 in_51_6
port 2 nsew signal input
rlabel m2 s 85 63 86 66 5 in_52_6
port 3 nsew signal input
rlabel m2 s 82 63 85 66 5 in_52_6
port 3 nsew signal input
rlabel m2 s 81 63 82 66 5 in_52_6
port 3 nsew signal input
rlabel m2 s 81 62 86 63 1 in_52_6
port 3 nsew signal input
rlabel m2 s 81 66 86 67 5 in_52_6
port 3 nsew signal input
rlabel m1 s 85 63 87 66 5 in_52_6
port 3 nsew signal input
rlabel m1 s 82 63 85 66 5 in_52_6
port 3 nsew signal input
rlabel m1 s 80 61 87 63 1 in_52_6
port 3 nsew signal input
rlabel m1 s 80 63 82 66 5 in_52_6
port 3 nsew signal input
rlabel m1 s 80 66 87 68 5 in_52_6
port 3 nsew signal input
rlabel m2 s 81 7 82 10 1 in_53_6
port 4 nsew signal input
rlabel m2 s 78 7 81 10 1 in_53_6
port 4 nsew signal input
rlabel m1 s 81 7 83 10 1 in_53_6
port 4 nsew signal input
rlabel m1 s 78 7 81 10 1 in_53_6
port 4 nsew signal input
rlabel m2 s 86 46 89 49 1 out
port 6 nsew signal output
rlabel m2 s 85 45 90 46 1 out
port 6 nsew signal output
rlabel m2 s 85 46 86 48 1 out
port 6 nsew signal output
rlabel m2 s 29 48 86 49 1 out
port 6 nsew signal output
rlabel m2 s 29 51 30 53 1 out
port 6 nsew signal output
rlabel m2 s 19 47 20 49 1 out
port 6 nsew signal output
rlabel m2 s 19 49 90 50 1 out
port 6 nsew signal output
rlabel m2 s 33 50 34 53 1 out
port 6 nsew signal output
rlabel m2 s 16 47 19 50 1 out
port 6 nsew signal output
rlabel m2 s 30 50 33 53 1 out
port 6 nsew signal output
rlabel m2 s 29 53 34 54 1 out
port 6 nsew signal output
rlabel m2 s 15 46 20 47 1 out
port 6 nsew signal output
rlabel m2 s 15 47 16 50 1 out
port 6 nsew signal output
rlabel m2 s 15 50 30 51 1 out
port 6 nsew signal output
rlabel m1 s 86 24 89 27 1 out
port 6 nsew signal output
rlabel m1 s 86 27 89 37 1 out
port 6 nsew signal output
rlabel m1 s 86 37 89 40 1 out
port 6 nsew signal output
rlabel m1 s 86 40 89 46 1 out
port 6 nsew signal output
rlabel m1 s 86 46 89 49 1 out
port 6 nsew signal output
rlabel m1 s 33 50 35 53 1 out
port 6 nsew signal output
rlabel m1 s 86 22 89 24 1 out
port 6 nsew signal output
rlabel m1 s 30 50 33 53 1 out
port 6 nsew signal output
rlabel m1 s 28 48 35 50 1 out
port 6 nsew signal output
rlabel m1 s 28 50 30 53 1 out
port 6 nsew signal output
rlabel m1 s 28 53 35 55 1 out
port 6 nsew signal output
rlabel m1 s 16 22 19 24 1 out
port 6 nsew signal output
rlabel m1 s 16 24 19 27 1 out
port 6 nsew signal output
rlabel m1 s 16 27 19 47 1 out
port 6 nsew signal output
rlabel m1 s 16 47 19 50 1 out
port 6 nsew signal output
rlabel m2 s 109 41 114 42 1 Vdd
port 2 nsew power input
rlabel m2 s 59 34 60 37 1 Vdd
port 2 nsew power input
rlabel m2 s 56 34 59 37 1 Vdd
port 2 nsew power input
rlabel m2 s 55 33 60 34 1 Vdd
port 2 nsew power input
rlabel m2 s 55 34 56 37 1 Vdd
port 2 nsew power input
rlabel m2 s 113 38 114 41 7 Vdd
port 2 nsew power input
rlabel m2 s 110 38 113 41 1 Vdd
port 2 nsew power input
rlabel m2 s 26 38 110 39 1 Vdd
port 2 nsew power input
rlabel m2 s 26 39 27 41 1 Vdd
port 2 nsew power input
rlabel m2 s 23 38 26 41 1 Vdd
port 2 nsew power input
rlabel m2 s 22 37 114 38 1 Vdd
port 2 nsew power input
rlabel m2 s 22 38 23 41 1 Vdd
port 2 nsew power input
rlabel m2 s 22 41 27 42 1 Vdd
port 2 nsew power input
rlabel m1 s 110 36 113 38 1 Vdd
port 2 nsew power input
rlabel m1 s 110 38 113 41 1 Vdd
port 2 nsew power input
rlabel m1 s 110 41 113 43 1 Vdd
port 2 nsew power input
rlabel m1 s 59 34 61 37 1 Vdd
port 2 nsew power input
rlabel m1 s 56 34 59 37 1 Vdd
port 2 nsew power input
rlabel m1 s 54 32 61 34 1 Vdd
port 2 nsew power input
rlabel m1 s 54 34 56 37 1 Vdd
port 2 nsew power input
rlabel m1 s 54 37 61 39 1 Vdd
port 2 nsew power input
rlabel m1 s 23 36 26 38 1 Vdd
port 2 nsew power input
rlabel m1 s 23 38 26 41 1 Vdd
port 2 nsew power input
rlabel m1 s 23 41 26 43 1 Vdd
port 2 nsew power input
rlabel m2 s 101 29 104 32 1 GND
port 1 nsew ground input
rlabel m2 s 100 28 105 29 1 GND
port 1 nsew ground input
rlabel m2 s 100 29 101 32 1 GND
port 1 nsew ground input
rlabel m2 s 100 32 105 33 1 GND
port 1 nsew ground input
rlabel m2 s 100 18 102 28 1 GND
port 1 nsew ground input
rlabel m2 s 74 14 75 16 1 GND
port 1 nsew ground input
rlabel m2 s 74 16 102 17 1 GND
port 1 nsew ground input
rlabel m2 s 71 14 74 17 1 GND
port 1 nsew ground input
rlabel m2 s 70 13 75 14 1 GND
port 1 nsew ground input
rlabel m2 s 70 14 71 16 1 GND
port 1 nsew ground input
rlabel m2 s 26 17 102 18 1 GND
port 1 nsew ground input
rlabel m2 s 26 18 27 20 1 GND
port 1 nsew ground input
rlabel m2 s 23 17 26 20 1 GND
port 1 nsew ground input
rlabel m2 s 22 16 71 17 1 GND
port 1 nsew ground input
rlabel m2 s 22 17 23 20 1 GND
port 1 nsew ground input
rlabel m2 s 22 20 27 21 1 GND
port 1 nsew ground input
rlabel m1 s 104 29 106 32 1 GND
port 1 nsew ground input
rlabel m1 s 101 29 104 32 1 GND
port 1 nsew ground input
rlabel m1 s 99 27 106 29 1 GND
port 1 nsew ground input
rlabel m1 s 99 29 101 32 1 GND
port 1 nsew ground input
rlabel m1 s 99 32 106 34 1 GND
port 1 nsew ground input
rlabel m1 s 71 26 74 28 1 GND
port 1 nsew ground input
rlabel m1 s 71 23 74 26 1 GND
port 1 nsew ground input
rlabel m1 s 23 26 26 28 1 GND
port 1 nsew ground input
rlabel m1 s 71 17 74 23 1 GND
port 1 nsew ground input
rlabel m1 s 71 14 74 17 1 GND
port 1 nsew ground input
rlabel m1 s 23 23 26 26 1 GND
port 1 nsew ground input
rlabel m1 s 23 17 26 20 1 GND
port 1 nsew ground input
rlabel m1 s 23 20 26 23 1 GND
port 1 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 120 72
string LEFclass CORE
string LEFsite CoreSite
string LEFsymmetry X Y
<< end >>
