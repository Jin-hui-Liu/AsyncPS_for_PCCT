magic
tech sky130A
magscale 1 2
timestamp 1753379664
<< nwell >>
rect 75 555 945 1035
rect 75 375 1320 555
rect 1575 375 1845 1035
<< nmos >>
rect 300 75 330 300
rect 405 210 435 300
rect 510 210 570 300
rect 915 210 945 300
rect 990 210 1320 300
rect 1425 75 1455 300
rect 1695 75 1725 300
<< pmos >>
rect 195 420 225 990
rect 300 420 330 990
rect 405 420 435 990
rect 510 420 570 570
rect 810 420 840 990
rect 915 420 945 510
rect 990 420 1200 510
rect 1695 420 1725 990
<< ndiff >>
rect 225 210 300 300
rect 225 165 240 210
rect 285 165 300 210
rect 225 75 300 165
rect 330 270 405 300
rect 330 225 345 270
rect 390 225 405 270
rect 330 210 405 225
rect 435 285 510 300
rect 435 240 450 285
rect 495 240 510 285
rect 435 210 510 240
rect 570 285 645 300
rect 570 240 585 285
rect 630 240 645 285
rect 570 210 645 240
rect 840 285 915 300
rect 840 240 855 285
rect 900 240 915 285
rect 840 210 915 240
rect 945 210 990 300
rect 1320 285 1425 300
rect 1320 240 1350 285
rect 1395 240 1425 285
rect 1320 210 1425 240
rect 330 75 390 210
rect 1365 75 1425 210
rect 1455 270 1530 300
rect 1455 225 1470 270
rect 1515 225 1530 270
rect 1455 75 1530 225
rect 1620 210 1695 300
rect 1620 165 1635 210
rect 1680 165 1695 210
rect 1620 75 1695 165
rect 1725 270 1800 300
rect 1725 225 1740 270
rect 1785 225 1800 270
rect 1725 75 1800 225
<< pdiff >>
rect 120 960 195 990
rect 120 915 135 960
rect 180 915 195 960
rect 120 420 195 915
rect 225 420 300 990
rect 330 420 405 990
rect 435 570 495 990
rect 735 885 810 990
rect 735 840 750 885
rect 795 840 810 885
rect 435 495 510 570
rect 435 450 450 495
rect 495 450 510 495
rect 435 420 510 450
rect 570 480 645 570
rect 570 435 585 480
rect 630 435 645 480
rect 570 420 645 435
rect 735 420 810 840
rect 840 510 900 990
rect 1620 960 1695 990
rect 1620 915 1635 960
rect 1680 915 1695 960
rect 840 480 915 510
rect 840 435 855 480
rect 900 435 915 480
rect 840 420 915 435
rect 945 420 990 510
rect 1200 480 1275 510
rect 1200 435 1215 480
rect 1260 435 1275 480
rect 1200 420 1275 435
rect 1620 420 1695 915
rect 1725 885 1800 990
rect 1725 840 1740 885
rect 1785 840 1800 885
rect 1725 420 1800 840
<< ndiffc >>
rect 240 165 285 210
rect 345 225 390 270
rect 450 240 495 285
rect 585 240 630 285
rect 855 240 900 285
rect 1350 240 1395 285
rect 1470 225 1515 270
rect 1635 165 1680 210
rect 1740 225 1785 270
<< pdiffc >>
rect 135 915 180 960
rect 750 840 795 885
rect 450 450 495 495
rect 585 435 630 480
rect 1635 915 1680 960
rect 855 435 900 480
rect 1215 435 1260 480
rect 1740 840 1785 885
<< poly >>
rect 270 1155 375 1185
rect 90 1110 195 1140
rect 90 1065 120 1110
rect 165 1065 195 1110
rect 270 1110 300 1155
rect 345 1110 375 1155
rect 270 1080 375 1110
rect 435 1095 540 1125
rect 90 1035 225 1065
rect 195 990 225 1035
rect 300 990 330 1080
rect 435 1050 465 1095
rect 510 1050 540 1095
rect 405 1020 540 1050
rect 765 1095 870 1125
rect 765 1050 795 1095
rect 840 1050 870 1095
rect 765 1020 870 1050
rect 1650 1110 1755 1140
rect 1650 1065 1680 1110
rect 1725 1065 1755 1110
rect 1650 1035 1755 1065
rect 405 990 435 1020
rect 810 990 840 1020
rect 1695 990 1725 1035
rect 510 570 570 600
rect 915 660 1035 690
rect 915 615 960 660
rect 1005 615 1035 660
rect 915 585 1035 615
rect 1080 615 1185 645
rect 915 510 945 585
rect 1080 570 1110 615
rect 1155 570 1185 615
rect 1080 540 1185 570
rect 990 510 1200 540
rect 195 390 225 420
rect 300 390 330 420
rect 300 300 330 330
rect 405 300 435 420
rect 510 300 570 420
rect 810 390 840 420
rect 915 300 945 420
rect 990 390 1200 420
rect 990 300 1320 330
rect 1425 300 1455 330
rect 1695 300 1725 420
rect 405 180 435 210
rect 510 120 570 210
rect 915 180 945 210
rect 990 180 1320 210
rect 1200 150 1305 180
rect 510 90 615 120
rect 300 15 330 75
rect 510 45 540 90
rect 585 45 615 90
rect 1200 105 1230 150
rect 1275 105 1305 150
rect 1200 75 1305 105
rect 1425 45 1455 75
rect 1695 45 1725 75
rect 510 15 615 45
rect 1395 15 1500 45
rect 225 -15 330 15
rect 225 -60 255 -15
rect 300 -60 330 -15
rect 1395 -30 1425 15
rect 1470 -30 1500 15
rect 1395 -60 1500 -30
rect 225 -90 330 -60
<< polycont >>
rect 120 1065 165 1110
rect 300 1110 345 1155
rect 465 1050 510 1095
rect 795 1050 840 1095
rect 1680 1065 1725 1110
rect 960 615 1005 660
rect 1110 570 1155 615
rect 540 45 585 90
rect 1230 105 1275 150
rect 255 -60 300 -15
rect 1425 -30 1470 15
<< locali >>
rect 270 1155 375 1185
rect 90 1110 195 1140
rect 90 1065 120 1110
rect 165 1065 195 1110
rect 270 1110 300 1155
rect 345 1110 375 1155
rect 270 1080 375 1110
rect 435 1095 540 1125
rect 90 1035 195 1065
rect 435 1050 465 1095
rect 510 1050 540 1095
rect 435 1020 540 1050
rect 765 1095 870 1125
rect 765 1050 795 1095
rect 840 1050 870 1095
rect 765 1020 870 1050
rect 1650 1110 1755 1140
rect 1650 1065 1680 1110
rect 1725 1065 1755 1110
rect 1650 1035 1755 1065
rect 135 960 180 990
rect 1635 960 1680 990
rect 135 885 180 915
rect 750 885 795 915
rect 1635 885 1680 915
rect 1740 885 1785 915
rect 750 810 795 840
rect 1740 810 1785 840
rect 930 660 1035 690
rect 930 615 960 660
rect 1005 615 1035 660
rect 930 585 1035 615
rect 1080 615 1185 645
rect 450 495 495 525
rect 450 420 495 450
rect 585 480 630 585
rect 1080 570 1110 615
rect 1155 570 1185 615
rect 1080 540 1185 570
rect 345 270 390 300
rect 240 210 285 240
rect 240 135 285 165
rect 345 105 390 225
rect 450 285 495 315
rect 450 210 495 240
rect 585 285 630 435
rect 585 210 630 240
rect 855 480 900 510
rect 855 285 900 435
rect 1095 330 1140 540
rect 1215 480 1260 510
rect 855 210 900 240
rect 1215 180 1260 435
rect 1350 285 1395 315
rect 1350 210 1395 240
rect 1470 270 1515 300
rect 1740 270 1785 300
rect 1470 195 1515 225
rect 1635 210 1680 240
rect 1200 150 1305 180
rect 510 90 615 120
rect 510 45 540 90
rect 585 45 615 90
rect 1200 105 1230 150
rect 1275 105 1305 150
rect 1740 195 1785 225
rect 1635 135 1680 165
rect 1200 75 1305 105
rect 510 15 615 45
rect 1395 15 1500 45
rect 225 -15 330 15
rect 225 -60 255 -15
rect 300 -60 330 -15
rect 1395 -30 1425 15
rect 1470 -30 1500 15
rect 1395 -60 1500 -30
rect 225 -90 330 -60
<< viali >>
rect 120 1065 165 1110
rect 300 1110 345 1155
rect 465 1050 510 1095
rect 795 1050 840 1095
rect 1680 1065 1725 1110
rect 135 915 180 960
rect 1635 915 1680 960
rect 750 840 795 885
rect 1740 840 1785 885
rect 585 585 630 630
rect 960 615 1005 660
rect 450 450 495 495
rect 240 165 285 210
rect 450 240 495 285
rect 1095 285 1140 330
rect 1215 435 1260 480
rect 1350 240 1395 285
rect 1470 225 1515 270
rect 345 60 390 105
rect 540 45 585 90
rect 1635 165 1680 210
rect 1740 225 1785 270
rect 255 -60 300 -15
rect 1425 -30 1470 15
<< metal1 >>
rect 285 1155 360 1170
rect 105 1110 180 1125
rect 105 1065 120 1110
rect 165 1065 180 1110
rect 285 1110 300 1155
rect 345 1110 360 1155
rect 1665 1110 1740 1125
rect 285 1095 360 1110
rect 450 1095 525 1110
rect 105 1050 180 1065
rect 450 1050 465 1095
rect 510 1050 525 1095
rect 450 1035 525 1050
rect 780 1095 855 1110
rect 780 1050 795 1095
rect 840 1050 855 1095
rect 1665 1065 1680 1110
rect 1725 1065 1740 1110
rect 1665 1050 1740 1065
rect 780 1035 855 1050
rect 120 960 1695 975
rect 120 915 135 960
rect 180 945 1635 960
rect 180 915 195 945
rect 120 900 195 915
rect 1620 915 1635 945
rect 1680 915 1695 960
rect 1620 900 1695 915
rect 735 885 810 900
rect 735 840 750 885
rect 795 855 810 885
rect 1725 885 1800 900
rect 1725 855 1740 885
rect 795 840 1740 855
rect 1785 840 1800 885
rect 735 825 1800 840
rect 945 660 1020 675
rect 945 645 960 660
rect 570 630 960 645
rect 570 585 585 630
rect 630 615 960 630
rect 1005 615 1020 660
rect 630 585 645 615
rect 945 600 1020 615
rect 570 570 645 585
rect 435 495 510 510
rect 435 450 450 495
rect 495 465 510 495
rect 1200 480 1275 495
rect 1200 465 1215 480
rect 495 450 1215 465
rect 435 435 1215 450
rect 1260 435 1275 480
rect 1200 420 1275 435
rect 1080 330 1155 345
rect 1080 300 1095 330
rect 435 285 1095 300
rect 1140 300 1155 330
rect 1140 285 1410 300
rect 435 240 450 285
rect 495 270 1350 285
rect 495 240 510 270
rect 435 225 510 240
rect 1335 240 1350 270
rect 1395 240 1410 285
rect 1335 225 1410 240
rect 1455 270 1800 285
rect 1455 225 1470 270
rect 1515 255 1740 270
rect 1515 225 1530 255
rect 1725 225 1740 255
rect 1785 225 1800 270
rect 225 210 300 225
rect 1455 210 1530 225
rect 1620 210 1695 225
rect 1725 210 1800 225
rect 225 165 240 210
rect 285 180 300 210
rect 1620 180 1635 210
rect 285 165 1635 180
rect 1680 165 1695 210
rect 225 150 1695 165
rect 330 105 405 120
rect 330 60 345 105
rect 390 75 405 105
rect 525 90 600 105
rect 525 75 540 90
rect 390 60 540 75
rect 330 45 540 60
rect 585 45 600 90
rect 525 30 600 45
rect 1410 15 1485 30
rect 240 -15 315 0
rect 240 -60 255 -15
rect 300 -60 315 -15
rect 1410 -30 1425 15
rect 1470 -30 1485 15
rect 1410 -45 1485 -30
rect 240 -75 315 -60
<< labels >>
flabel ndiff 270 75 270 75 1 FreeSerif 120 0 0 0 #4
flabel ndiff 375 75 375 75 1 FreeSerif 120 0 0 0 out
flabel ndiff 1365 210 1365 210 1 FreeSerif 120 0 0 0 GND
flabel ndiff 1500 75 1500 75 1 FreeSerif 120 0 0 0 #5
flabel ndiff 1770 75 1770 75 1 FreeSerif 120 0 0 0 #5
flabel ndiff 1665 75 1665 75 1 FreeSerif 120 0 0 0 #4
flabel poly 1695 345 1695 345 3 FreeSerif 120 0 0 0 in(3)
flabel poly 1425 315 1425 315 3 FreeSerif 120 0 0 0 in(5)
flabel poly 1005 315 1005 315 3 FreeSerif 120 0 0 0 Vdd
flabel poly 1005 405 1005 405 3 FreeSerif 120 0 0 0 GND
flabel poly 915 360 915 360 3 FreeSerif 120 0 0 0 #16
flabel poly 810 405 810 405 3 FreeSerif 120 0 0 0 in(4)
flabel poly 510 360 510 360 3 FreeSerif 120 0 0 0 out
flabel poly 405 360 405 360 3 FreeSerif 120 0 0 0 in(0)
flabel poly 300 405 300 405 3 FreeSerif 120 0 0 0 in(1)
flabel poly 300 315 300 315 3 FreeSerif 120 0 0 0 in(6)
flabel poly 195 405 195 405 3 FreeSerif 120 0 0 0 in(2)
flabel ndiff 480 210 480 210 1 FreeSerif 120 0 0 0 GND
flabel ndiff 615 210 615 210 1 FreeSerif 120 0 0 0 #16
flabel ndiff 885 210 885 210 1 FreeSerif 120 0 0 0 out
flabel pdiff 1770 420 1770 420 1 FreeSerif 120 0 0 0 #9
flabel pdiff 1665 420 1665 420 1 FreeSerif 120 0 0 0 #10
flabel pdiff 1245 420 1245 420 1 FreeSerif 120 0 0 0 Vdd
flabel pdiff 885 420 885 420 1 FreeSerif 120 0 0 0 out
flabel pdiff 780 420 780 420 1 FreeSerif 120 0 0 0 #9
flabel pdiff 615 420 615 420 1 FreeSerif 120 0 0 0 #16
flabel pdiff 480 420 480 420 1 FreeSerif 120 0 0 0 Vdd
flabel pdiff 165 420 165 420 1 FreeSerif 120 0 0 0 #10
flabel metal1 1125 330 1125 330 1 FreeSerif 120 0 0 0 GND
port 1 n
flabel metal1 1260 495 1260 495 1 FreeSerif 120 0 0 0 Vdd
port 2 n
flabel metal1 270 -75 270 -75 5 FreeSerif 120 0 0 0 in(6)
port 3 s
flabel metal1 1455 -45 1455 -45 5 FreeSerif 120 0 0 0 in(5)
port 4 s
flabel metal1 825 1110 825 1110 1 FreeSerif 120 0 0 0 in(4)
port 5 n
flabel metal1 1710 1125 1710 1125 1 FreeSerif 120 0 0 0 in(3)
port 6 n
flabel metal1 135 1125 135 1125 1 FreeSerif 120 0 0 0 in(2)
port 7 n
flabel metal1 315 1170 315 1170 1 FreeSerif 120 0 0 0 in(1)
port 8 n
flabel metal1 570 30 570 30 5 FreeSerif 120 0 0 0 out
port 9 s
flabel metal1 495 1110 495 1110 1 FreeSerif 120 0 0 0 in(0)
port 10 n
<< end >>
