magic
tech sky130l
timestamp 1753821931
<< checkpaint >>

<< nwell >>

<< labels >>

<< end >>
