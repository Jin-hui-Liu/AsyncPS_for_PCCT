magic
tech sky130A
magscale 1 2
timestamp 1753015926
<< checkpaint >>
rect -1140 1725 2640 2040
rect -1140 1695 2895 1725
rect -1140 -915 2970 1695
rect -1140 -945 2895 -915
rect -1140 -1110 2715 -945
rect -1140 -1140 2640 -1110
rect -1140 -1170 2595 -1140
rect -1140 -1200 2535 -1170
<< nmos >>
rect 300 150 330 240
rect 405 150 465 240
rect 705 150 1035 240
rect 1140 90 1170 240
rect 1245 90 1275 240
rect 1350 150 1380 240
<< pmos >>
rect 195 345 225 690
rect 300 345 330 690
rect 405 345 465 495
rect 1245 345 1275 690
rect 1350 345 1380 435
rect 1425 345 1635 435
<< ndiff >>
rect 225 150 300 240
rect 330 150 405 240
rect 465 150 540 240
rect 630 150 705 240
rect 1035 150 1140 240
rect 1080 90 1140 150
rect 1170 90 1245 240
rect 1275 150 1350 240
rect 1380 150 1455 240
rect 1275 90 1335 150
<< pdiff >>
rect 120 345 195 690
rect 225 345 300 690
rect 330 495 390 690
rect 330 345 405 495
rect 465 345 540 495
rect 1170 345 1245 690
rect 1275 435 1335 690
rect 1275 345 1350 435
rect 1380 345 1425 435
rect 1635 345 1710 435
<< poly >>
rect 195 690 225 720
rect 300 690 330 720
rect 1245 690 1275 720
rect 405 495 465 525
rect 1350 435 1380 465
rect 1425 435 1635 465
rect 195 315 225 345
rect 300 315 330 345
rect 405 315 465 345
rect 1245 315 1275 345
rect 1350 315 1380 345
rect 1425 315 1635 345
rect 300 240 330 270
rect 405 240 465 270
rect 705 240 1035 270
rect 1140 240 1170 270
rect 1245 240 1275 270
rect 1350 240 1380 270
rect 300 120 330 150
rect 405 120 465 150
rect 705 120 1035 150
rect 1350 120 1380 150
rect 1140 60 1170 90
rect 1245 60 1275 90
<< metal1 >>
rect 120 720 180 780
rect 360 720 420 780
rect 600 720 660 780
rect 840 720 900 780
rect 1080 720 1140 780
rect 1320 720 1380 780
rect 120 60 180 120
<< labels >>
rlabel pdiff 467 347 467 347 3 #10
rlabel ndiff 467 152 467 152 3 #10
rlabel poly 407 242 407 242 3 out
rlabel poly 407 317 407 317 3 out
rlabel ndiff 332 152 332 152 3 GND
rlabel pdiff 332 347 332 347 3 Vdd
rlabel poly 302 242 302 242 3 in(0)
rlabel poly 302 317 302 317 3 in(0)
rlabel ndiff 227 152 227 152 3 out
rlabel poly 197 317 197 317 3 in(1)
rlabel pdiff 122 347 122 347 3 #7
rlabel pdiff 1637 347 1637 347 3 Vdd
rlabel poly 1427 317 1427 317 3 GND
rlabel ndiff 1382 152 1382 152 3 #12
rlabel poly 1352 242 1352 242 3 #10
rlabel poly 1352 317 1352 317 3 #10
rlabel pdiff 1277 347 1277 347 3 out
rlabel ndiff 1277 92 1277 92 3 out
rlabel poly 1247 242 1247 242 3 in(2)
rlabel poly 1247 317 1247 317 3 in(2)
rlabel pdiff 1172 347 1172 347 3 #7
rlabel poly 1142 242 1142 242 3 in(3)
rlabel ndiff 1037 152 1037 152 3 GND
rlabel poly 707 242 707 242 3 Vdd
rlabel ndiff 632 152 632 152 3 #12
rlabel metal1 1322 722 1322 722 3 GND
port 1 e
rlabel metal1 1082 722 1082 722 3 Vdd
port 2 e
rlabel metal1 842 722 842 722 3 in(3)
port 3 e
rlabel metal1 602 722 602 722 3 in(2)
port 4 e
rlabel metal1 362 722 362 722 3 in(1)
port 5 e
rlabel metal1 122 62 122 62 3 out
port 6 e
rlabel metal1 122 722 122 722 3 in(0)
port 7 e
<< end >>
