magic
tech sky130A
timestamp 1753015928
<< checkpaint >>
rect 57870 555120 509130 567630
rect 57870 510120 509130 531630
rect 57870 426870 509130 459630
rect 57870 321120 509130 362880
rect 57870 226620 509130 257130
rect 57870 127620 509130 169380
rect 57870 39870 509130 63630
<< nwell >>
rect 58500 555750 508500 567000
rect 58500 510750 508500 531000
rect 58500 427500 508500 459000
rect 58500 321750 508500 362250
rect 58500 227250 508500 256500
rect 58500 128250 508500 168750
rect 58500 40500 508500 63000
<< labels >>
rlabel nwell 58501 40501 58501 40501 3 Vdd
rlabel nwell 58501 128251 58501 128251 3 Vdd
rlabel nwell 58501 227251 58501 227251 3 Vdd
rlabel nwell 58501 321751 58501 321751 3 Vdd
rlabel nwell 58501 427501 58501 427501 3 Vdd
rlabel nwell 58501 510751 58501 510751 3 Vdd
rlabel nwell 58501 555751 58501 555751 3 Vdd
<< end >>
