VERSION 5.6 ;

BUSBITCHARS "[]" ;

DIVIDERCHAR "/" ;

UNITS
    DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005000 ; 

CLEARANCEMEASURE EUCLIDEAN ; 

USEMINSPACING OBS ON ; 

SITE CoreSite
    CLASS CORE ;
    SIZE 0.600000 BY 0.300000 ;
END CoreSite

LAYER li
   TYPE ROUTING ;
   DIRECTION VERTICAL ;
   MINWIDTH 0.300000 ;
   AREA 0.056250 ;
   WIDTH 0.300000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 0.225000 ;
   PITCH 0.600000 0.600000 ;
END li

LAYER mcon
    TYPE CUT ;
    SPACING 0.225000 ;
    WIDTH 0.300000 ;
    ENCLOSURE ABOVE 0.075000 0.075000 ;
    ENCLOSURE BELOW 0.000000 0.000000 ;
END mcon

LAYER met1
   TYPE ROUTING ;
   DIRECTION HORIZONTAL ;
   MINWIDTH 0.150000 ;
   AREA 0.084375 ;
   WIDTH 0.150000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 0.150000 ;
   PITCH 0.300000 0.300000 ;
END met1

LAYER v1
    TYPE CUT ;
    SPACING 0.075000 ;
    WIDTH 0.300000 ;
    ENCLOSURE ABOVE 0.075000 0.075000 ;
    ENCLOSURE BELOW 0.075000 0.075000 ;
END v1

LAYER met2
   TYPE ROUTING ;
   DIRECTION VERTICAL ;
   MINWIDTH 0.150000 ;
   AREA 0.073125 ;
   WIDTH 0.150000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 0.150000 ;
   PITCH 0.300000 0.300000 ;
END met2

LAYER v2
    TYPE CUT ;
    SPACING 0.150000 ;
    WIDTH 0.300000 ;
    ENCLOSURE ABOVE 0.075000 0.075000 ;
    ENCLOSURE BELOW 0.075000 0.000000 ;
END v2

LAYER met3
   TYPE ROUTING ;
   DIRECTION HORIZONTAL ;
   MINWIDTH 0.300000 ;
   AREA 0.241875 ;
   WIDTH 0.300000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 0.300000 ;
   PITCH 0.600000 0.600000 ;
END met3

LAYER v3
    TYPE CUT ;
    SPACING 0.150000 ;
    WIDTH 0.450000 ;
    ENCLOSURE ABOVE 0.075000 0.075000 ;
    ENCLOSURE BELOW 0.075000 0.000000 ;
END v3

LAYER met4
   TYPE ROUTING ;
   DIRECTION VERTICAL ;
   MINWIDTH 0.300000 ;
   AREA 0.241875 ;
   WIDTH 0.300000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 0.300000 ;
   PITCH 0.600000 0.600000 ;
END met4

LAYER v4
    TYPE CUT ;
    SPACING 0.450000 ;
    WIDTH 1.200000 ;
    ENCLOSURE ABOVE 0.150000 0.150000 ;
    ENCLOSURE BELOW 0.000000 0.000000 ;
END v4

LAYER met5
   TYPE ROUTING ;
   DIRECTION HORIZONTAL ;
   MINWIDTH 1.650000 ;
   AREA 4.005000 ;
   WIDTH 1.650000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 1.650000 ;
   PITCH 3.300000 3.300000 ;
END met5

LAYER OVERLAP
   TYPE OVERLAP ;
END OVERLAP

VIA mcon_C DEFAULT
   LAYER li ;
     RECT -0.150000 -0.150000 0.150000 0.150000 ;
   LAYER mcon ;
     RECT -0.150000 -0.150000 0.150000 0.150000 ;
   LAYER met1 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END mcon_C

VIA v1_C DEFAULT
   LAYER met1 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v1 ;
     RECT -0.150000 -0.150000 0.150000 0.150000 ;
   LAYER met2 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v1_C

VIA v2_C DEFAULT
   LAYER met2 ;
     RECT -0.150000 -0.225000 0.150000 0.225000 ;
   LAYER v2 ;
     RECT -0.150000 -0.150000 0.150000 0.150000 ;
   LAYER met3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v2_C

VIA v2_Ch
   LAYER met2 ;
     RECT -0.225000 -0.150000 0.225000 0.150000 ;
   LAYER v2 ;
     RECT -0.150000 -0.150000 0.150000 0.150000 ;
   LAYER met3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v2_Ch

VIA v2_Cv
   LAYER met2 ;
     RECT -0.150000 -0.225000 0.150000 0.225000 ;
   LAYER v2 ;
     RECT -0.150000 -0.150000 0.150000 0.150000 ;
   LAYER met3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v2_Cv

VIA v3_C DEFAULT
   LAYER met3 ;
     RECT -0.300000 -0.225000 0.300000 0.225000 ;
   LAYER v3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER met4 ;
     RECT -0.300000 -0.300000 0.300000 0.300000 ;
END v3_C

VIA v3_Ch
   LAYER met3 ;
     RECT -0.300000 -0.225000 0.300000 0.225000 ;
   LAYER v3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER met4 ;
     RECT -0.300000 -0.300000 0.300000 0.300000 ;
END v3_Ch

VIA v3_Cv
   LAYER met3 ;
     RECT -0.300000 -0.225000 0.300000 0.225000 ;
   LAYER v3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER met4 ;
     RECT -0.300000 -0.300000 0.300000 0.300000 ;
END v3_Cv

VIA v4_C DEFAULT
   LAYER met4 ;
     RECT -0.600000 -0.600000 0.600000 0.600000 ;
   LAYER v4 ;
     RECT -0.600000 -0.600000 0.600000 0.600000 ;
   LAYER met5 ;
     RECT -0.750000 -0.750000 0.750000 0.750000 ;
END v4_C

MACRO _0_0cell_0_0ginvx0
    CLASS CORE ;
    FOREIGN _0_0cell_0_0ginvx0 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.400000 BY 2.700000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN in_50_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 0.600000 2.100000 0.900000 2.400000 ;
        END
    END in_50_6
    PIN out
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 0.600000 0.300000 0.900000 0.600000 ;
        END
        ANTENNADIFFAREA 0.393750 ;
    END out
    PIN Vdd
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER li ;
        RECT 1.200000 2.100000 1.500000 2.400000 ;
        END
        ANTENNADIFFAREA 0.225000 ;
    END Vdd
    PIN GND
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER li ;
        RECT 1.800000 2.100000 2.100000 2.400000 ;
        END
        ANTENNADIFFAREA 0.168750 ;
    END GND
END _0_0cell_0_0ginvx0

MACRO _0_0cell_0_0g0n1n2n3naaa_04256aaaox0
    CLASS CORE ;
    FOREIGN _0_0cell_0_0g0n1n2n3naaa_04256aaaox0 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 9.600000 BY 5.400000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN in_50_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 0.600000 4.800000 0.900000 5.100000 ;
        END
    END in_50_6
    PIN in_51_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 1.200000 4.800000 1.500000 5.100000 ;
        END
    END in_51_6
    PIN in_52_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 1.800000 4.800000 2.100000 5.100000 ;
        END
    END in_52_6
    PIN in_53_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 2.400000 4.800000 2.700000 5.100000 ;
        END
    END in_53_6
    PIN in_54_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 3.000000 4.800000 3.300000 5.100000 ;
        END
    END in_54_6
    PIN in_55_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 3.600000 4.800000 3.900000 5.100000 ;
        END
    END in_55_6
    PIN in_56_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 4.200000 4.800000 4.500000 5.100000 ;
        END
    END in_56_6
    PIN out
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 0.600000 0.300000 0.900000 0.600000 ;
        END
        ANTENNADIFFAREA 1.293750 ;
    END out
    PIN Vdd
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER li ;
        RECT 4.800000 4.800000 5.100000 5.100000 ;
        END
        ANTENNADIFFAREA 0.843750 ;
    END Vdd
    PIN GND
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER li ;
        RECT 5.400000 4.800000 5.700000 5.100000 ;
        END
        ANTENNADIFFAREA 0.270000 ;
    END GND
    OBS
      LAYER li ;
         RECT 0.600000 1.800000 8.925000 3.525000 ;
    END
END _0_0cell_0_0g0n1n2n3naaa_04256aaaox0

MACRO _0_0cell_0_0g0n1n2n3n4naaao_025a4267aaooax0
    CLASS CORE ;
    FOREIGN _0_0cell_0_0g0n1n2n3n4naaao_025a4267aaooax0 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 12.600000 BY 6.000000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN in_50_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 0.600000 5.400000 0.900000 5.700000 ;
        END
    END in_50_6
    PIN in_51_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 1.800000 5.400000 2.100000 5.700000 ;
        END
    END in_51_6
    PIN in_52_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 3.000000 5.400000 3.300000 5.700000 ;
        END
    END in_52_6
    PIN in_53_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 4.200000 5.400000 4.500000 5.700000 ;
        END
    END in_53_6
    PIN in_54_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 5.400000 5.400000 5.700000 5.700000 ;
        END
    END in_54_6
    PIN in_55_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 6.600000 5.400000 6.900000 5.700000 ;
        END
    END in_55_6
    PIN in_56_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 7.800000 5.400000 8.100000 5.700000 ;
        END
    END in_56_6
    PIN in_57_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 9.000000 5.400000 9.300000 5.700000 ;
        END
    END in_57_6
    PIN out
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 0.600000 0.300000 0.900000 0.600000 ;
        END
        ANTENNADIFFAREA 2.182500 ;
    END out
    PIN Vdd
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER li ;
        RECT 10.200000 5.400000 10.500000 5.700000 ;
        END
        ANTENNADIFFAREA 0.236250 ;
    END Vdd
    PIN GND
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER li ;
        RECT 11.400000 5.400000 11.700000 5.700000 ;
        END
        ANTENNADIFFAREA 0.618750 ;
    END GND
    OBS
      LAYER li ;
         RECT 0.600000 1.800000 11.925000 4.125000 ;
    END
END _0_0cell_0_0g0n1n2n3n4naaao_025a4267aaooax0

MACRO _0_0cell_0_0g0n1n2n3naaa_02ox0
    CLASS CORE ;
    FOREIGN _0_0cell_0_0g0n1n2n3naaa_02ox0 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 9.000000 BY 4.500000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN in_50_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 0.600000 3.900000 0.900000 4.200000 ;
        END
    END in_50_6
    PIN in_51_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 1.800000 3.900000 2.100000 4.200000 ;
        END
    END in_51_6
    PIN in_52_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 3.000000 3.900000 3.300000 4.200000 ;
        END
    END in_52_6
    PIN in_53_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 4.200000 3.900000 4.500000 4.200000 ;
        END
    END in_53_6
    PIN out
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 0.600000 0.300000 0.900000 0.600000 ;
        END
        ANTENNADIFFAREA 1.518750 ;
    END out
    PIN Vdd
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER li ;
        RECT 5.400000 3.900000 5.700000 4.200000 ;
        END
        ANTENNADIFFAREA 0.843750 ;
    END Vdd
    PIN GND
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER li ;
        RECT 6.600000 3.900000 6.900000 4.200000 ;
        END
        ANTENNADIFFAREA 0.337500 ;
    END GND
    OBS
      LAYER li ;
         RECT 0.600000 1.800000 8.325000 2.625000 ;
    END
END _0_0cell_0_0g0n1n2n3naaa_02ox0

MACRO _0_0cell_0_0g0n1n2n3n4n5naaaaa_0653aaox0
    CLASS CORE ;
    FOREIGN _0_0cell_0_0g0n1n2n3n4n5naaaaa_0653aaox0 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 10.800000 BY 6.000000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN in_50_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 0.600000 5.400000 0.900000 5.700000 ;
        END
    END in_50_6
    PIN in_51_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 1.800000 5.400000 2.100000 5.700000 ;
        END
    END in_51_6
    PIN in_52_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 3.000000 5.400000 3.300000 5.700000 ;
        END
    END in_52_6
    PIN in_53_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 4.200000 5.400000 4.500000 5.700000 ;
        END
    END in_53_6
    PIN in_54_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 5.400000 5.400000 5.700000 5.700000 ;
        END
    END in_54_6
    PIN in_55_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 6.600000 5.400000 6.900000 5.700000 ;
        END
    END in_55_6
    PIN in_56_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 7.800000 5.400000 8.100000 5.700000 ;
        END
    END in_56_6
    PIN out
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 0.600000 0.300000 0.900000 0.600000 ;
        END
        ANTENNADIFFAREA 2.193750 ;
    END out
    PIN Vdd
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER li ;
        RECT 9.000000 5.400000 9.300000 5.700000 ;
        END
        ANTENNADIFFAREA 1.181250 ;
    END Vdd
    PIN GND
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER li ;
        RECT 10.200000 5.400000 10.500000 5.700000 ;
        END
        ANTENNADIFFAREA 0.270000 ;
    END GND
    OBS
      LAYER li ;
         RECT 0.600000 1.800000 10.125000 4.125000 ;
    END
END _0_0cell_0_0g0n1n2n3n4n5naaaaa_0653aaox0

MACRO _0_0cell_0_0g0n1n2n3n4naaaa_0536aaox0
    CLASS CORE ;
    FOREIGN _0_0cell_0_0g0n1n2n3n4naaaa_0536aaox0 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 9.600000 BY 5.700000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN in_50_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 0.600000 5.100000 0.900000 5.400000 ;
        END
    END in_50_6
    PIN in_51_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 1.200000 5.100000 1.500000 5.400000 ;
        END
    END in_51_6
    PIN in_52_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 1.800000 5.100000 2.100000 5.400000 ;
        END
    END in_52_6
    PIN in_53_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 2.400000 5.100000 2.700000 5.400000 ;
        END
    END in_53_6
    PIN in_54_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 3.000000 5.100000 3.300000 5.400000 ;
        END
    END in_54_6
    PIN in_55_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 3.600000 5.100000 3.900000 5.400000 ;
        END
    END in_55_6
    PIN in_56_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 4.200000 5.100000 4.500000 5.400000 ;
        END
    END in_56_6
    PIN out
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 0.600000 0.300000 0.900000 0.600000 ;
        END
        ANTENNADIFFAREA 1.361250 ;
    END out
    PIN Vdd
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER li ;
        RECT 4.800000 5.100000 5.100000 5.400000 ;
        END
        ANTENNADIFFAREA 1.023750 ;
    END Vdd
    PIN GND
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER li ;
        RECT 5.400000 5.100000 5.700000 5.400000 ;
        END
        ANTENNADIFFAREA 0.270000 ;
    END GND
    OBS
      LAYER li ;
         RECT 0.600000 1.800000 8.925000 3.825000 ;
    END
END _0_0cell_0_0g0n1n2n3n4naaaa_0536aaox0

MACRO _0_0cell_0_0ginvx1
    CLASS CORE ;
    FOREIGN _0_0cell_0_0ginvx1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 2.400000 BY 3.000000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN in_50_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 0.600000 2.400000 0.900000 2.700000 ;
        END
    END in_50_6
    PIN out
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 0.600000 0.300000 0.900000 0.600000 ;
        END
        ANTENNADIFFAREA 0.450000 ;
    END out
    PIN Vdd
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER li ;
        RECT 1.200000 2.400000 1.500000 2.700000 ;
        END
        ANTENNADIFFAREA 0.281250 ;
    END Vdd
    PIN GND
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER li ;
        RECT 1.800000 2.400000 2.100000 2.700000 ;
        END
        ANTENNADIFFAREA 0.168750 ;
    END GND
END _0_0cell_0_0ginvx1

MACRO _0_0cell_0_0g0n1n2naa_032aox0
    CLASS CORE ;
    FOREIGN _0_0cell_0_0g0n1n2naa_032aox0 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 9.000000 BY 4.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN in_50_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 0.600000 3.600000 0.900000 3.900000 ;
        END
    END in_50_6
    PIN in_51_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 1.800000 3.600000 2.100000 3.900000 ;
        END
    END in_51_6
    PIN in_52_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 3.000000 3.600000 3.300000 3.900000 ;
        END
    END in_52_6
    PIN in_53_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 4.200000 3.600000 4.500000 3.900000 ;
        END
    END in_53_6
    PIN out
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 0.600000 0.300000 0.900000 0.600000 ;
        END
        ANTENNADIFFAREA 0.911250 ;
    END out
    PIN Vdd
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER li ;
        RECT 5.400000 3.600000 5.700000 3.900000 ;
        END
        ANTENNADIFFAREA 0.686250 ;
    END Vdd
    PIN GND
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER li ;
        RECT 6.600000 3.600000 6.900000 3.900000 ;
        END
        ANTENNADIFFAREA 0.270000 ;
    END GND
    OBS
      LAYER li ;
         RECT 0.600000 1.800000 8.325000 2.325000 ;
    END
END _0_0cell_0_0g0n1n2naa_032aox0

MACRO _0_0cell_0_0g0n1n2na3n2n4n5naaa2n6n7naaooa_082a92aoox0
    CLASS CORE ;
    FOREIGN _0_0cell_0_0g0n1n2na3n2n4n5naaa2n6n7naaooa_082a92aoox0 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 12.600000 BY 6.000000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN in_50_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 0.600000 5.400000 0.900000 5.700000 ;
        END
    END in_50_6
    PIN in_51_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 1.200000 5.400000 1.500000 5.700000 ;
        END
    END in_51_6
    PIN in_52_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 1.800000 5.400000 2.100000 5.700000 ;
        END
    END in_52_6
    PIN in_53_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 2.400000 5.400000 2.700000 5.700000 ;
        END
    END in_53_6
    PIN in_54_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 3.000000 5.400000 3.300000 5.700000 ;
        END
    END in_54_6
    PIN in_55_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 3.600000 5.400000 3.900000 5.700000 ;
        END
    END in_55_6
    PIN in_56_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 4.200000 5.400000 4.500000 5.700000 ;
        END
    END in_56_6
    PIN in_57_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 4.800000 5.400000 5.100000 5.700000 ;
        END
    END in_57_6
    PIN in_58_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 5.400000 5.400000 5.700000 5.700000 ;
        END
    END in_58_6
    PIN in_59_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 6.000000 5.400000 6.300000 5.700000 ;
        END
    END in_59_6
    PIN out
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 0.600000 0.300000 0.900000 0.600000 ;
        END
        ANTENNADIFFAREA 2.137500 ;
    END out
    PIN Vdd
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER li ;
        RECT 6.600000 5.400000 6.900000 5.700000 ;
        END
        ANTENNADIFFAREA 1.023750 ;
    END Vdd
    PIN GND
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER li ;
        RECT 7.200000 5.400000 7.500000 5.700000 ;
        END
        ANTENNADIFFAREA 0.551250 ;
    END GND
    OBS
      LAYER li ;
         RECT 0.600000 1.800000 11.925000 4.125000 ;
    END
END _0_0cell_0_0g0n1n2na3n2n4n5naaa2n6n7naaooa_082a92aoox0

MACRO welltap_svt
    CLASS CORE WELLTAP ;
    FOREIGN welltap_svt 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.200000 BY 2.100000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Vdd
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER li ;
        RECT 0.600000 1.500000 0.900000 1.800000 ;
        END
    END Vdd
    PIN GND
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER li ;
        RECT 0.600000 0.300000 0.900000 0.600000 ;
        END
    END GND
END welltap_svt

MACRO circuitppnp
   CLASS CORE ;
   FOREIGN circuitppnp 0.000000 0.000000 ;
   ORIGIN 0.000000 0.000000 ; 
   SIZE 65.400000 BY 70.200000 ; 
   SYMMETRY X Y ;
   SITE CoreSite ;
END circuitppnp

MACRO circuitwell
   CLASS CORE ;
   FOREIGN circuitwell 0.000000 0.000000 ;
   ORIGIN 0.000000 0.000000 ; 
   SIZE 65.400000 BY 70.200000 ; 
   SYMMETRY X Y ;
   SITE CoreSite ;
END circuitwell

