magic
tech sky130A
magscale 1 2
timestamp 1753299154
<< nwell >>
rect 75 435 1260 795
rect 75 255 1740 435
<< nmos >>
rect 300 90 330 180
rect 405 90 465 180
rect 705 90 1035 180
rect 1110 90 1140 180
rect 1380 90 1410 180
<< pmos >>
rect 195 300 225 750
rect 300 300 330 750
rect 405 300 465 450
rect 705 300 735 750
rect 1110 300 1140 750
rect 1380 300 1410 390
rect 1455 300 1620 390
<< ndiff >>
rect 225 165 300 180
rect 225 120 240 165
rect 285 120 300 165
rect 225 90 300 120
rect 330 165 405 180
rect 330 120 345 165
rect 390 120 405 165
rect 330 90 405 120
rect 465 165 540 180
rect 465 120 480 165
rect 525 120 540 165
rect 465 90 540 120
rect 630 165 705 180
rect 630 120 645 165
rect 690 120 705 165
rect 630 90 705 120
rect 1035 165 1110 180
rect 1035 120 1050 165
rect 1095 120 1110 165
rect 1035 90 1110 120
rect 1140 165 1215 180
rect 1140 120 1155 165
rect 1200 120 1215 165
rect 1140 90 1215 120
rect 1305 165 1380 180
rect 1305 120 1320 165
rect 1365 120 1380 165
rect 1305 90 1380 120
rect 1410 165 1485 180
rect 1410 120 1425 165
rect 1470 120 1485 165
rect 1410 90 1485 120
<< pdiff >>
rect 120 705 195 750
rect 120 660 135 705
rect 180 660 195 705
rect 120 300 195 660
rect 225 300 300 750
rect 330 450 390 750
rect 630 555 705 750
rect 630 510 645 555
rect 690 510 705 555
rect 330 375 405 450
rect 330 330 345 375
rect 390 330 405 375
rect 330 300 405 330
rect 465 360 540 450
rect 465 315 480 360
rect 525 315 540 360
rect 465 300 540 315
rect 630 300 705 510
rect 735 300 1110 750
rect 1140 705 1215 750
rect 1140 660 1155 705
rect 1200 660 1215 705
rect 1140 300 1215 660
rect 1305 360 1380 390
rect 1305 315 1320 360
rect 1365 315 1380 360
rect 1305 300 1380 315
rect 1410 300 1455 390
rect 1620 375 1695 390
rect 1620 330 1635 375
rect 1680 330 1695 375
rect 1620 300 1695 330
<< ndiffc >>
rect 240 120 285 165
rect 345 120 390 165
rect 480 120 525 165
rect 645 120 690 165
rect 1050 120 1095 165
rect 1155 120 1200 165
rect 1320 120 1365 165
rect 1425 120 1470 165
<< pdiffc >>
rect 135 660 180 705
rect 645 510 690 555
rect 345 330 390 375
rect 480 315 525 360
rect 1155 660 1200 705
rect 1320 315 1365 360
rect 1635 330 1680 375
<< poly >>
rect 120 855 225 885
rect 120 810 150 855
rect 195 810 225 855
rect 120 780 225 810
rect 195 750 225 780
rect 300 855 405 885
rect 300 810 330 855
rect 375 810 405 855
rect 300 780 405 810
rect 630 855 735 885
rect 630 810 660 855
rect 705 810 735 855
rect 630 780 735 810
rect 300 750 330 780
rect 705 750 735 780
rect 1110 855 1215 885
rect 1110 810 1140 855
rect 1185 810 1215 855
rect 1110 780 1215 810
rect 1110 750 1140 780
rect 420 555 525 585
rect 420 510 450 555
rect 495 510 525 555
rect 420 480 525 510
rect 405 450 465 480
rect 1380 390 1410 420
rect 1455 390 1620 420
rect 195 270 225 300
rect 300 180 330 300
rect 405 180 465 300
rect 705 270 735 300
rect 705 180 1035 210
rect 1110 180 1140 300
rect 1380 180 1410 300
rect 1455 270 1620 300
rect 1515 225 1620 270
rect 1515 180 1545 225
rect 1590 180 1620 225
rect 1515 150 1620 180
rect 300 60 330 90
rect 405 60 465 90
rect 705 60 1035 90
rect 1110 60 1140 90
rect 825 30 930 60
rect 1380 45 1410 90
rect 825 -15 855 30
rect 900 -15 930 30
rect 825 -45 930 -15
rect 1305 15 1410 45
rect 1305 -30 1335 15
rect 1380 -30 1410 15
rect 1305 -60 1410 -30
<< polycont >>
rect 150 810 195 855
rect 330 810 375 855
rect 660 810 705 855
rect 1140 810 1185 855
rect 450 510 495 555
rect 1545 180 1590 225
rect 855 -15 900 30
rect 1335 -30 1380 15
<< locali >>
rect 120 855 225 885
rect 120 810 150 855
rect 195 810 225 855
rect 120 780 225 810
rect 300 855 405 885
rect 300 810 330 855
rect 375 810 405 855
rect 300 780 405 810
rect 630 855 735 885
rect 630 810 660 855
rect 705 810 735 855
rect 630 780 735 810
rect 1110 855 1215 885
rect 1110 810 1140 855
rect 1185 810 1215 855
rect 1110 780 1215 810
rect 135 705 180 735
rect 135 630 180 660
rect 1155 705 1200 735
rect 1155 630 1200 660
rect 420 555 525 585
rect 420 510 450 555
rect 495 510 525 555
rect 420 480 525 510
rect 645 555 690 585
rect 645 480 690 510
rect 240 165 285 465
rect 345 375 390 405
rect 345 300 390 330
rect 480 360 525 390
rect 240 90 285 120
rect 345 165 390 195
rect 345 90 390 120
rect 480 165 525 315
rect 480 60 525 120
rect 645 165 690 195
rect 645 90 690 120
rect 855 60 900 345
rect 1050 165 1095 195
rect 1050 90 1095 120
rect 1155 165 1200 510
rect 1155 90 1200 120
rect 1320 360 1365 510
rect 1320 165 1365 315
rect 1635 375 1680 405
rect 1635 300 1680 330
rect 1515 225 1620 255
rect 1320 90 1365 120
rect 1425 165 1470 195
rect 1515 180 1545 225
rect 1590 180 1620 225
rect 1515 150 1620 180
rect 1425 90 1470 120
rect 480 0 525 15
rect 825 30 930 60
rect 825 -15 855 30
rect 900 -15 930 30
rect 825 -45 930 -15
rect 1305 15 1410 45
rect 1305 -30 1335 15
rect 1380 -30 1410 15
rect 1305 -60 1410 -30
<< viali >>
rect 150 810 195 855
rect 330 810 375 855
rect 660 810 705 855
rect 1140 810 1185 855
rect 135 660 180 705
rect 1155 660 1200 705
rect 450 510 495 555
rect 240 465 285 510
rect 645 510 690 555
rect 1155 510 1200 555
rect 345 330 390 375
rect 345 195 390 240
rect 855 345 900 390
rect 645 120 690 165
rect 1050 195 1095 240
rect 1320 510 1365 555
rect 1635 330 1680 375
rect 1425 120 1470 165
rect 1545 180 1590 225
rect 480 15 525 60
rect 1335 -30 1380 15
<< metal1 >>
rect 135 855 210 870
rect 135 810 150 855
rect 195 810 210 855
rect 135 795 210 810
rect 315 855 390 870
rect 315 810 330 855
rect 375 810 390 855
rect 315 795 390 810
rect 645 855 720 870
rect 645 810 660 855
rect 705 810 720 855
rect 645 795 720 810
rect 1125 855 1200 870
rect 1125 810 1140 855
rect 1185 810 1200 855
rect 1125 795 1200 810
rect 120 705 1215 720
rect 120 660 135 705
rect 180 690 1155 705
rect 180 660 195 690
rect 120 645 195 660
rect 1140 660 1155 690
rect 1200 660 1215 705
rect 1140 645 1215 660
rect 435 555 510 570
rect 435 525 450 555
rect 225 510 450 525
rect 495 525 510 555
rect 630 555 705 570
rect 630 525 645 555
rect 495 510 645 525
rect 690 525 705 555
rect 1140 555 1215 570
rect 1140 525 1155 555
rect 690 510 1155 525
rect 1200 525 1215 555
rect 1305 555 1380 570
rect 1305 525 1320 555
rect 1200 510 1320 525
rect 1365 510 1380 555
rect 225 465 240 510
rect 285 495 1380 510
rect 285 465 300 495
rect 225 450 300 465
rect 840 390 915 405
rect 330 375 405 390
rect 840 375 855 390
rect 330 330 345 375
rect 390 345 855 375
rect 900 375 915 390
rect 1620 375 1695 390
rect 900 345 1635 375
rect 390 330 405 345
rect 840 330 915 345
rect 1620 330 1635 345
rect 1680 330 1695 375
rect 330 315 405 330
rect 1620 315 1695 330
rect 330 240 1605 255
rect 330 195 345 240
rect 390 225 1050 240
rect 390 195 405 225
rect 330 180 405 195
rect 1035 195 1050 225
rect 1095 225 1605 240
rect 1095 195 1110 225
rect 1515 210 1545 225
rect 1035 180 1110 195
rect 1530 180 1545 210
rect 1590 180 1605 225
rect 630 165 705 180
rect 630 120 645 165
rect 690 135 705 165
rect 1410 165 1485 180
rect 1530 165 1605 180
rect 1410 135 1425 165
rect 690 120 1425 135
rect 1470 120 1485 165
rect 630 105 1485 120
rect 465 60 540 75
rect 465 15 480 60
rect 525 30 540 60
rect 525 15 1395 30
rect 465 0 1335 15
rect 1320 -30 1335 0
rect 1380 -30 1395 15
rect 1320 -45 1395 -30
<< labels >>
flabel poly 1380 240 1380 240 3 FreeSerif 120 0 0 0 #10
flabel poly 1470 285 1470 285 3 FreeSerif 120 0 0 0 GND
flabel pdiff 1635 300 1635 300 1 FreeSerif 120 0 0 0 Vdd
flabel ndiff 1455 90 1455 90 1 FreeSerif 120 0 0 0 #12
flabel ndiff 1350 90 1350 90 1 FreeSerif 120 0 0 0 out
flabel ndiff 1185 90 1185 90 1 FreeSerif 120 0 0 0 out
flabel ndiff 1080 90 1080 90 1 FreeSerif 120 0 0 0 GND
flabel poly 735 195 735 195 1 FreeSerif 120 0 0 0 Vdd
flabel ndiff 675 90 675 90 1 FreeSerif 120 0 0 0 #12
flabel ndiff 510 90 510 90 1 FreeSerif 120 0 0 0 #10
flabel ndiff 375 90 375 90 1 FreeSerif 120 0 0 0 GND
flabel ndiff 270 90 270 90 1 FreeSerif 120 0 0 0 out
flabel poly 195 285 195 285 3 FreeSerif 120 0 0 0 in(1)
flabel poly 300 240 300 240 3 FreeSerif 120 0 0 0 in(0)
flabel poly 405 240 405 240 3 FreeSerif 120 0 0 0 out
flabel poly 705 285 705 285 3 FreeSerif 120 0 0 0 in(3)
flabel pdiff 675 300 675 300 1 FreeSerif 120 0 0 0 out
flabel pdiff 375 300 375 300 1 FreeSerif 120 0 0 0 Vdd
flabel pdiff 165 300 165 300 1 FreeSerif 120 0 0 0 #6
flabel pdiff 510 300 510 300 1 FreeSerif 120 0 0 0 #10
flabel pdiff 1185 300 1185 300 1 FreeSerif 120 0 0 0 #6
flabel pdiff 1350 300 1350 300 1 FreeSerif 120 0 0 0 out
flabel poly 1110 240 1110 240 3 FreeSerif 120 0 0 0 in(2)
flabel metal1 1605 210 1605 210 3 FreeSerif 120 0 0 0 GND
port 1 e
flabel metal1 885 405 885 405 1 FreeSerif 120 0 0 0 Vdd
port 2 n
flabel metal1 675 870 675 870 1 FreeSerif 120 0 0 0 in(3)
port 3 n
flabel metal1 1170 870 1170 870 1 FreeSerif 120 0 0 0 in(2)
port 4 n
flabel metal1 165 870 165 870 1 FreeSerif 120 0 0 0 in(1)
port 5 n
flabel metal1 480 570 480 570 1 FreeSerif 120 0 0 0 out
port 6 n
flabel metal1 360 870 360 870 1 FreeSerif 120 0 0 0 in(0)
port 7 n
<< end >>
