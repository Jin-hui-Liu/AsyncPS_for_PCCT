magic
tech sky130A
magscale 1 2
timestamp 1753015926
<< checkpaint >>
rect -1140 1740 3600 2400
rect -1140 -870 3675 1740
rect -1140 -900 3600 -870
rect -1140 -1080 3030 -900
rect -1140 -1110 2955 -1080
rect -1140 -1185 1785 -1110
rect -1140 -1200 1725 -1185
rect -930 -1215 1725 -1200
<< nmos >>
rect 195 285 225 480
rect 330 75 360 480
rect 435 75 465 480
rect 540 375 570 480
rect 675 180 705 480
rect 810 390 870 480
rect 1530 330 1560 480
rect 1665 180 1695 480
rect 1935 390 1965 480
rect 2010 390 2340 480
<< pmos >>
rect 435 585 465 1035
rect 540 585 570 1035
rect 675 585 705 705
rect 810 585 870 735
rect 1110 585 1320 675
rect 1425 585 1455 1035
rect 1530 585 1560 1035
rect 1935 585 1965 675
<< ndiff >>
rect 120 285 195 480
rect 225 285 330 480
rect 270 75 330 285
rect 360 75 435 480
rect 465 375 540 480
rect 570 375 675 480
rect 465 75 525 375
rect 615 180 675 375
rect 705 390 810 480
rect 870 390 945 480
rect 705 180 765 390
rect 1455 330 1530 480
rect 1560 330 1665 480
rect 1605 180 1665 330
rect 1695 180 1770 480
rect 1860 390 1935 480
rect 1965 390 2010 480
rect 2340 390 2415 480
<< pdiff >>
rect 360 585 435 1035
rect 465 585 540 1035
rect 570 705 630 1035
rect 750 705 810 735
rect 570 585 675 705
rect 705 585 810 705
rect 870 585 945 735
rect 1365 675 1425 1035
rect 1035 585 1110 675
rect 1320 585 1425 675
rect 1455 585 1530 1035
rect 1560 585 1635 1035
rect 1860 585 1935 675
rect 1965 585 2040 675
<< poly >>
rect 435 1035 465 1065
rect 540 1035 570 1065
rect 1425 1035 1455 1065
rect 1530 1035 1560 1065
rect 810 735 870 765
rect 675 705 705 735
rect 1110 675 1320 705
rect 1935 675 1965 705
rect 435 555 465 585
rect 540 555 570 585
rect 675 555 705 585
rect 810 555 870 585
rect 1110 555 1320 585
rect 1425 555 1455 585
rect 1530 555 1560 585
rect 1935 555 1965 585
rect 195 480 225 510
rect 330 480 360 510
rect 435 480 465 510
rect 540 480 570 510
rect 675 480 705 510
rect 810 480 870 510
rect 1530 480 1560 510
rect 1665 480 1695 510
rect 1935 480 1965 510
rect 2010 480 2340 510
rect 195 255 225 285
rect 540 345 570 375
rect 810 360 870 390
rect 1530 300 1560 330
rect 1935 360 1965 390
rect 2010 360 2340 390
rect 675 150 705 180
rect 1665 150 1695 180
rect 330 45 360 75
rect 435 45 465 75
<< metal1 >>
rect 120 1080 180 1140
rect 360 1080 420 1140
rect 600 1080 660 1140
rect 840 1080 900 1140
rect 1080 1080 1140 1140
rect 1320 1080 1380 1140
rect 1560 1080 1620 1140
rect 1800 1080 1860 1140
rect 2040 1080 2100 1140
rect 2280 1080 2340 1140
rect 120 60 180 120
<< labels >>
rlabel poly 812 482 812 482 3 out
rlabel poly 812 557 812 557 3 out
rlabel pdiff 872 587 872 587 3 #18
rlabel ndiff 872 392 872 392 3 #18
rlabel poly 677 482 677 482 3 in(0)
rlabel poly 677 557 677 557 3 in(0)
rlabel pdiff 707 587 707 587 3 Vdd
rlabel ndiff 707 182 707 182 3 GND
rlabel ndiff 572 377 572 377 3 #3
rlabel poly 542 482 542 482 3 in(4)
rlabel poly 542 557 542 557 3 in(4)
rlabel pdiff 572 587 572 587 3 out
rlabel ndiff 467 77 467 77 3 out
rlabel poly 437 482 437 482 3 in(7)
rlabel poly 437 557 437 557 3 in(3)
rlabel pdiff 362 587 362 587 3 #14
rlabel poly 332 482 332 482 3 in(6)
rlabel poly 197 482 197 482 3 in(2)
rlabel ndiff 122 287 122 287 3 #3
rlabel pdiff 1562 587 1562 587 3 #14
rlabel ndiff 1697 182 1697 182 3 out
rlabel poly 1667 482 1667 482 3 in(5)
rlabel poly 1532 557 1532 557 3 in(2)
rlabel poly 1532 482 1532 482 3 in(2)
rlabel poly 1427 557 1427 557 3 in(1)
rlabel ndiff 1457 332 1457 332 3 #3
rlabel pdiff 1322 587 1322 587 3 Vdd
rlabel poly 1112 557 1112 557 3 GND
rlabel pdiff 1037 587 1037 587 3 #19
rlabel ndiff 2342 392 2342 392 3 GND
rlabel poly 2012 482 2012 482 3 Vdd
rlabel pdiff 1967 587 1967 587 3 out
rlabel poly 1937 482 1937 482 3 #18
rlabel poly 1937 557 1937 557 3 #18
rlabel ndiff 1862 392 1862 392 3 out
rlabel pdiff 1862 587 1862 587 3 #19
rlabel metal1 2282 1082 2282 1082 3 GND
port 1 e
rlabel metal1 2042 1082 2042 1082 3 Vdd
port 2 e
rlabel metal1 1802 1082 1802 1082 3 in(7)
port 3 e
rlabel metal1 1562 1082 1562 1082 3 in(6)
port 4 e
rlabel metal1 1322 1082 1322 1082 3 in(5)
port 5 e
rlabel metal1 1082 1082 1082 1082 3 in(4)
port 6 e
rlabel metal1 842 1082 842 1082 3 in(3)
port 7 e
rlabel metal1 602 1082 602 1082 3 in(2)
port 8 e
rlabel metal1 362 1082 362 1082 3 in(1)
port 9 e
rlabel metal1 122 62 122 62 3 out
port 10 e
rlabel metal1 122 1082 122 1082 3 in(0)
port 11 e
<< end >>
