magic
tech sky130A
magscale 1 2
timestamp 1753015926
<< checkpaint >>
rect -1140 -180 3360 2400
rect -1140 -1185 3300 -180
rect -1140 -1200 3225 -1185
rect 30 -1215 3225 -1200
<< nmos >>
rect 375 210 405 300
rect 480 210 540 300
rect 780 210 810 300
rect 855 210 1185 300
rect 1290 75 1320 300
rect 1665 75 1695 300
rect 1935 75 1965 300
<< pmos >>
rect 195 405 225 1080
rect 270 405 300 1080
rect 375 405 405 1080
rect 480 405 540 555
rect 780 405 810 495
rect 855 405 1065 495
rect 1560 405 1590 1080
rect 1665 405 1695 1080
rect 1935 405 1965 1080
<< ndiff >>
rect 300 210 375 300
rect 405 210 480 300
rect 540 210 615 300
rect 705 210 780 300
rect 810 210 855 300
rect 1185 210 1290 300
rect 1230 75 1290 210
rect 1320 75 1395 300
rect 1590 75 1665 300
rect 1695 75 1770 300
rect 1860 75 1935 300
rect 1965 75 2040 300
<< pdiff >>
rect 120 405 195 1080
rect 225 405 270 1080
rect 300 405 375 1080
rect 405 555 465 1080
rect 405 405 480 555
rect 540 405 615 555
rect 705 405 780 495
rect 810 405 855 495
rect 1065 405 1140 495
rect 1485 405 1560 1080
rect 1590 405 1665 1080
rect 1695 405 1770 1080
rect 1860 405 1935 1080
rect 1965 405 2040 1080
<< poly >>
rect 195 1080 225 1110
rect 270 1080 300 1110
rect 375 1080 405 1110
rect 1560 1080 1590 1110
rect 1665 1080 1695 1110
rect 1935 1080 1965 1110
rect 480 555 540 585
rect 780 495 810 525
rect 855 495 1065 525
rect 195 375 225 405
rect 270 375 300 405
rect 375 375 405 405
rect 480 375 540 405
rect 780 375 810 405
rect 855 375 1065 405
rect 1560 375 1590 405
rect 1665 375 1695 405
rect 1935 375 1965 405
rect 375 300 405 330
rect 480 300 540 330
rect 780 300 810 330
rect 855 300 1185 330
rect 1290 300 1320 330
rect 1665 300 1695 330
rect 1935 300 1965 330
rect 375 180 405 210
rect 480 180 540 210
rect 780 180 810 210
rect 855 180 1185 210
rect 1290 45 1320 75
rect 1665 45 1695 75
rect 1935 45 1965 75
<< metal1 >>
rect 120 1080 180 1140
rect 360 1080 420 1140
rect 600 1080 660 1140
rect 840 1080 900 1140
rect 1080 1080 1140 1140
rect 1320 1080 1380 1140
rect 1560 1080 1620 1140
rect 1800 1080 1860 1140
rect 2040 1080 2100 1140
rect 120 60 180 120
<< labels >>
rlabel pdiff 542 407 542 407 3 #17
rlabel poly 482 377 482 377 3 out
rlabel ndiff 542 212 542 212 3 #17
rlabel pdiff 407 407 407 407 3 Vdd
rlabel poly 482 302 482 302 3 out
rlabel poly 377 377 377 377 3 in(0)
rlabel ndiff 407 212 407 212 3 GND
rlabel poly 377 302 377 302 3 in(0)
rlabel poly 272 377 272 377 3 in(1)
rlabel ndiff 302 212 302 212 3 out
rlabel poly 197 377 197 377 3 in(2)
rlabel pdiff 122 407 122 407 3 #11
rlabel poly 1292 302 1292 302 3 in(6)
rlabel ndiff 1322 77 1322 77 3 #5
rlabel ndiff 1187 212 1187 212 3 GND
rlabel pdiff 1067 407 1067 407 3 Vdd
rlabel poly 857 302 857 302 3 Vdd
rlabel poly 857 377 857 377 3 GND
rlabel poly 782 302 782 302 3 #17
rlabel poly 782 377 782 377 3 #17
rlabel ndiff 707 212 707 212 3 out
rlabel pdiff 707 407 707 407 3 out
rlabel ndiff 1697 77 1697 77 3 #4
rlabel pdiff 1697 407 1697 407 3 #11
rlabel poly 1667 302 1667 302 3 in(3)
rlabel poly 1667 377 1667 377 3 in(3)
rlabel ndiff 1592 77 1592 77 3 out
rlabel poly 1562 377 1562 377 3 in(4)
rlabel pdiff 1487 407 1487 407 3 #9
rlabel ndiff 1967 77 1967 77 3 #5
rlabel pdiff 1967 407 1967 407 3 #9
rlabel poly 1937 302 1937 302 3 in(5)
rlabel poly 1937 377 1937 377 3 in(5)
rlabel ndiff 1862 77 1862 77 3 #4
rlabel pdiff 1862 407 1862 407 3 out
rlabel metal1 2042 1082 2042 1082 3 GND
port 1 e
rlabel metal1 1802 1082 1802 1082 3 Vdd
port 2 e
rlabel metal1 1562 1082 1562 1082 3 in(6)
port 3 e
rlabel metal1 1322 1082 1322 1082 3 in(5)
port 4 e
rlabel metal1 1082 1082 1082 1082 3 in(4)
port 5 e
rlabel metal1 842 1082 842 1082 3 in(3)
port 6 e
rlabel metal1 602 1082 602 1082 3 in(2)
port 7 e
rlabel metal1 362 1082 362 1082 3 in(1)
port 8 e
rlabel metal1 122 62 122 62 3 out
port 9 e
rlabel metal1 122 1082 122 1082 3 in(0)
port 10 e
<< end >>
