magic
tech sky130l
timestamp 1753821931
<< m1 >>
rect 550 991 554 1008
rect 128 911 132 955
rect 128 803 132 907
rect 472 895 476 907
rect 168 787 172 799
rect 168 763 172 783
rect 512 755 516 767
rect 512 751 536 755
rect 640 747 644 783
rect 800 739 804 815
rect 848 755 852 779
rect 856 747 860 759
rect 264 687 268 691
rect 256 683 268 687
rect 256 639 260 683
rect 328 643 332 663
rect 168 567 172 583
rect 256 571 260 635
rect 472 635 476 663
rect 824 643 828 711
rect 1012 694 1016 719
rect 80 535 84 542
rect 168 535 172 563
rect 296 555 300 571
rect 168 511 172 531
rect 392 531 396 563
rect 496 455 500 563
rect 520 511 524 571
rect 552 495 556 583
rect 792 543 796 583
rect 152 395 156 447
rect 1012 382 1016 399
rect 408 291 412 323
rect 448 211 452 267
rect 136 179 140 199
rect 456 191 460 243
rect 592 163 596 203
rect 632 155 636 167
rect 484 143 492 147
rect 488 139 492 143
rect 632 143 636 151
rect 488 135 496 139
rect 552 99 556 131
rect 550 95 556 99
rect 550 72 554 95
<< m2c >>
rect 111 989 115 993
rect 550 987 554 991
rect 959 989 963 993
rect 111 971 115 975
rect 959 971 963 975
rect 128 955 132 959
rect 111 909 115 913
rect 128 907 132 911
rect 111 891 115 895
rect 111 829 115 833
rect 111 811 115 815
rect 472 907 476 911
rect 959 909 963 913
rect 472 891 476 895
rect 959 891 963 895
rect 959 829 963 833
rect 800 815 804 819
rect 128 799 132 803
rect 168 799 172 803
rect 168 783 172 787
rect 640 783 644 787
rect 168 759 172 763
rect 512 767 516 771
rect 536 751 540 755
rect 640 743 644 747
rect 959 811 963 815
rect 848 779 852 783
rect 848 751 852 755
rect 856 759 860 763
rect 856 743 860 747
rect 800 735 804 739
rect 1012 719 1016 723
rect 824 711 828 715
rect 111 705 115 709
rect 264 691 268 695
rect 111 687 115 691
rect 328 663 332 667
rect 328 639 332 643
rect 472 663 476 667
rect 256 635 260 639
rect 111 617 115 621
rect 111 599 115 603
rect 168 583 172 587
rect 959 705 963 709
rect 959 687 963 691
rect 824 639 828 643
rect 472 631 476 635
rect 959 617 963 621
rect 959 599 963 603
rect 552 583 556 587
rect 256 567 260 571
rect 296 571 300 575
rect 168 563 172 567
rect 80 531 84 535
rect 520 571 524 575
rect 296 551 300 555
rect 392 563 396 567
rect 168 531 172 535
rect 392 527 396 531
rect 496 563 500 567
rect 168 507 172 511
rect 111 485 115 489
rect 111 467 115 471
rect 520 507 524 511
rect 792 583 796 587
rect 792 539 796 543
rect 552 491 556 495
rect 959 485 963 489
rect 959 467 963 471
rect 496 451 500 455
rect 152 447 156 451
rect 111 405 115 409
rect 959 405 963 409
rect 152 391 156 395
rect 1012 399 1016 403
rect 111 387 115 391
rect 959 387 963 391
rect 408 323 412 327
rect 111 293 115 297
rect 959 293 963 297
rect 408 287 412 291
rect 111 275 115 279
rect 959 275 963 279
rect 448 267 452 271
rect 111 213 115 217
rect 448 207 452 211
rect 456 243 460 247
rect 136 199 140 203
rect 111 195 115 199
rect 959 213 963 217
rect 456 187 460 191
rect 592 203 596 207
rect 136 175 140 179
rect 959 195 963 199
rect 592 159 596 163
rect 632 167 636 171
rect 632 151 636 155
rect 480 143 484 147
rect 632 139 636 143
rect 496 135 500 139
rect 552 131 556 135
rect 111 117 115 121
rect 111 99 115 103
rect 959 117 963 121
rect 959 99 963 103
<< m2 >>
rect 134 1000 140 1001
rect 134 996 135 1000
rect 139 996 140 1000
rect 134 995 140 996
rect 318 1000 324 1001
rect 318 996 319 1000
rect 323 996 324 1000
rect 318 995 324 996
rect 526 1000 532 1001
rect 526 996 527 1000
rect 531 996 532 1000
rect 526 995 532 996
rect 734 1000 740 1001
rect 734 996 735 1000
rect 739 996 740 1000
rect 926 1000 932 1001
rect 926 996 927 1000
rect 931 996 932 1000
rect 734 995 740 996
rect 834 995 840 996
rect 926 995 932 996
rect 110 993 116 994
rect 110 989 111 993
rect 115 989 116 993
rect 110 988 116 989
rect 549 991 555 992
rect 549 987 550 991
rect 554 990 555 991
rect 834 991 835 995
rect 839 991 840 995
rect 834 990 840 991
rect 958 993 964 994
rect 554 988 838 990
rect 958 989 959 993
rect 963 989 964 993
rect 958 988 964 989
rect 554 987 555 988
rect 549 986 555 987
rect 938 987 944 988
rect 938 986 939 987
rect 744 984 939 986
rect 202 979 208 980
rect 744 979 746 984
rect 938 983 939 984
rect 943 983 944 987
rect 938 982 944 983
rect 946 979 952 980
rect 202 978 203 979
rect 145 976 203 978
rect 110 975 116 976
rect 110 971 111 975
rect 115 971 116 975
rect 202 975 203 976
rect 207 975 208 979
rect 946 978 947 979
rect 202 974 208 975
rect 232 976 329 978
rect 432 976 537 978
rect 937 976 947 978
rect 110 970 116 971
rect 134 968 140 969
rect 134 964 135 968
rect 139 964 140 968
rect 232 966 234 976
rect 149 964 234 966
rect 318 968 324 969
rect 318 964 319 968
rect 323 964 324 968
rect 432 966 434 976
rect 946 975 947 976
rect 951 975 952 979
rect 946 974 952 975
rect 958 975 964 976
rect 938 971 944 972
rect 333 964 434 966
rect 526 968 532 969
rect 526 964 527 968
rect 531 964 532 968
rect 734 968 740 969
rect 926 968 932 969
rect 134 963 140 964
rect 318 963 324 964
rect 526 963 532 964
rect 127 959 133 960
rect 127 955 128 959
rect 132 958 133 959
rect 426 959 432 960
rect 132 956 334 958
rect 132 955 133 956
rect 127 954 133 955
rect 286 951 292 952
rect 286 947 287 951
rect 291 947 292 951
rect 286 946 292 947
rect 298 951 304 952
rect 298 947 299 951
rect 303 947 304 951
rect 318 951 324 952
rect 318 950 319 951
rect 313 948 319 950
rect 298 946 304 947
rect 318 947 319 948
rect 323 947 324 951
rect 332 949 334 956
rect 426 955 427 959
rect 431 958 432 959
rect 536 958 538 965
rect 734 964 735 968
rect 739 964 740 968
rect 758 967 764 968
rect 758 966 759 967
rect 749 964 759 966
rect 734 963 740 964
rect 758 963 759 964
rect 763 963 764 967
rect 926 964 927 968
rect 931 964 932 968
rect 938 967 939 971
rect 943 967 944 971
rect 958 971 959 975
rect 963 971 964 975
rect 958 970 964 971
rect 938 966 944 967
rect 926 963 932 964
rect 758 962 764 963
rect 431 956 538 958
rect 431 955 432 956
rect 426 954 432 955
rect 442 951 448 952
rect 442 950 443 951
rect 393 948 443 950
rect 318 946 324 947
rect 442 947 443 948
rect 447 947 448 951
rect 442 946 448 947
rect 298 927 304 928
rect 298 926 299 927
rect 224 924 299 926
rect 134 920 140 921
rect 158 920 164 921
rect 182 920 188 921
rect 224 920 226 924
rect 298 923 299 924
rect 303 926 304 927
rect 303 924 734 926
rect 303 923 304 924
rect 298 922 304 923
rect 230 920 236 921
rect 454 920 460 921
rect 518 920 524 921
rect 582 920 588 921
rect 646 920 652 921
rect 710 920 716 921
rect 134 916 135 920
rect 139 916 140 920
rect 134 915 140 916
rect 146 919 152 920
rect 146 915 147 919
rect 151 915 152 919
rect 158 916 159 920
rect 163 916 164 920
rect 158 915 164 916
rect 170 919 176 920
rect 170 915 171 919
rect 175 915 176 919
rect 182 916 183 920
rect 187 916 188 920
rect 222 919 228 920
rect 222 918 223 919
rect 197 916 223 918
rect 182 915 188 916
rect 222 915 223 916
rect 227 915 228 919
rect 230 916 231 920
rect 235 916 236 920
rect 250 919 256 920
rect 250 918 251 919
rect 245 916 251 918
rect 230 915 236 916
rect 250 915 251 916
rect 255 918 256 919
rect 298 919 304 920
rect 298 918 299 919
rect 255 916 299 918
rect 255 915 256 916
rect 146 914 152 915
rect 170 914 176 915
rect 222 914 228 915
rect 250 914 256 915
rect 298 915 299 916
rect 303 915 304 919
rect 454 916 455 920
rect 459 916 460 920
rect 454 915 460 916
rect 466 919 472 920
rect 466 915 467 919
rect 471 915 472 919
rect 518 916 519 920
rect 523 916 524 920
rect 518 915 524 916
rect 530 919 536 920
rect 530 915 531 919
rect 535 915 536 919
rect 582 916 583 920
rect 587 916 588 920
rect 630 919 636 920
rect 630 918 631 919
rect 597 916 631 918
rect 582 915 588 916
rect 630 915 631 916
rect 635 915 636 919
rect 646 916 647 920
rect 651 916 652 920
rect 666 919 672 920
rect 666 918 667 919
rect 661 916 667 918
rect 646 915 652 916
rect 666 915 667 916
rect 671 915 672 919
rect 710 916 711 920
rect 715 916 716 920
rect 710 915 716 916
rect 722 919 728 920
rect 722 915 723 919
rect 727 915 728 919
rect 298 914 304 915
rect 466 914 472 915
rect 530 914 536 915
rect 630 914 636 915
rect 666 914 672 915
rect 722 914 728 915
rect 110 913 116 914
rect 110 909 111 913
rect 115 909 116 913
rect 310 912 316 913
rect 110 908 116 909
rect 127 911 133 912
rect 127 907 128 911
rect 132 910 133 911
rect 132 908 145 910
rect 310 908 311 912
rect 315 908 316 912
rect 132 907 133 908
rect 127 906 133 907
rect 190 907 196 908
rect 168 898 170 905
rect 190 903 191 907
rect 195 903 196 907
rect 190 902 196 903
rect 238 907 244 908
rect 310 907 316 908
rect 370 911 376 912
rect 370 907 371 911
rect 375 910 376 911
rect 471 911 477 912
rect 471 910 472 911
rect 375 908 472 910
rect 375 907 376 908
rect 238 903 239 907
rect 243 903 244 907
rect 370 906 376 907
rect 471 907 472 908
rect 476 907 477 911
rect 732 910 734 924
rect 766 920 772 921
rect 822 920 828 921
rect 886 920 892 921
rect 926 920 932 921
rect 766 916 767 920
rect 771 916 772 920
rect 814 919 820 920
rect 814 918 815 919
rect 781 916 815 918
rect 766 915 772 916
rect 814 915 815 916
rect 819 915 820 919
rect 822 916 823 920
rect 827 916 828 920
rect 822 915 828 916
rect 834 919 840 920
rect 834 915 835 919
rect 839 915 840 919
rect 886 916 887 920
rect 891 916 892 920
rect 918 919 924 920
rect 918 918 919 919
rect 901 916 919 918
rect 886 915 892 916
rect 918 915 919 916
rect 923 915 924 919
rect 926 916 927 920
rect 931 916 932 920
rect 946 919 952 920
rect 946 918 947 919
rect 941 916 947 918
rect 926 915 932 916
rect 946 915 947 916
rect 951 915 952 919
rect 814 914 820 915
rect 834 914 840 915
rect 918 914 924 915
rect 946 914 952 915
rect 958 913 964 914
rect 732 908 777 910
rect 958 909 959 913
rect 963 909 964 913
rect 958 908 964 909
rect 471 906 477 907
rect 538 907 544 908
rect 238 902 244 903
rect 378 903 384 904
rect 250 899 256 900
rect 250 898 251 899
rect 168 896 251 898
rect 110 895 116 896
rect 110 891 111 895
rect 115 891 116 895
rect 250 895 251 896
rect 255 895 256 899
rect 378 899 379 903
rect 383 902 384 903
rect 510 903 516 904
rect 510 902 511 903
rect 383 900 511 902
rect 383 899 384 900
rect 378 898 384 899
rect 510 899 511 900
rect 515 902 516 903
rect 528 902 530 905
rect 538 903 539 907
rect 543 906 544 907
rect 654 907 660 908
rect 543 904 593 906
rect 543 903 544 904
rect 538 902 544 903
rect 654 903 655 907
rect 659 903 660 907
rect 654 902 660 903
rect 702 907 708 908
rect 702 903 703 907
rect 707 906 708 907
rect 842 907 848 908
rect 842 906 843 907
rect 707 904 721 906
rect 833 904 843 906
rect 707 903 708 904
rect 702 902 708 903
rect 842 903 843 904
rect 847 903 848 907
rect 946 907 952 908
rect 946 906 947 907
rect 842 902 848 903
rect 515 900 530 902
rect 515 899 516 900
rect 510 898 516 899
rect 834 899 840 900
rect 250 894 256 895
rect 310 895 316 896
rect 110 890 116 891
rect 310 891 311 895
rect 315 891 316 895
rect 310 890 316 891
rect 471 895 477 896
rect 471 891 472 895
rect 476 894 477 895
rect 530 895 536 896
rect 530 894 531 895
rect 476 892 531 894
rect 476 891 477 892
rect 471 890 477 891
rect 530 891 531 892
rect 535 891 536 895
rect 834 895 835 899
rect 839 898 840 899
rect 896 898 898 905
rect 937 904 947 906
rect 946 903 947 904
rect 951 903 952 907
rect 946 902 952 903
rect 839 896 898 898
rect 839 895 840 896
rect 834 894 840 895
rect 958 895 964 896
rect 530 890 536 891
rect 958 891 959 895
rect 963 891 964 895
rect 958 890 964 891
rect 134 888 140 889
rect 134 884 135 888
rect 139 884 140 888
rect 134 883 140 884
rect 158 888 164 889
rect 158 884 159 888
rect 163 884 164 888
rect 158 883 164 884
rect 182 888 188 889
rect 182 884 183 888
rect 187 884 188 888
rect 182 883 188 884
rect 230 888 236 889
rect 230 884 231 888
rect 235 884 236 888
rect 458 888 464 889
rect 458 884 459 888
rect 463 884 464 888
rect 230 883 236 884
rect 426 883 432 884
rect 458 883 464 884
rect 518 888 524 889
rect 518 884 519 888
rect 523 884 524 888
rect 518 883 524 884
rect 582 888 588 889
rect 582 884 583 888
rect 587 884 588 888
rect 582 883 588 884
rect 646 888 652 889
rect 646 884 647 888
rect 651 884 652 888
rect 646 883 652 884
rect 710 888 716 889
rect 710 884 711 888
rect 715 884 716 888
rect 710 883 716 884
rect 766 888 772 889
rect 766 884 767 888
rect 771 884 772 888
rect 766 883 772 884
rect 822 888 828 889
rect 822 884 823 888
rect 827 884 828 888
rect 822 883 828 884
rect 886 888 892 889
rect 886 884 887 888
rect 891 884 892 888
rect 886 883 892 884
rect 926 888 932 889
rect 926 884 927 888
rect 931 884 932 888
rect 926 883 932 884
rect 426 882 427 883
rect 317 880 427 882
rect 126 879 132 880
rect 126 875 127 879
rect 131 878 132 879
rect 190 879 196 880
rect 190 878 191 879
rect 131 876 191 878
rect 131 875 132 876
rect 126 874 132 875
rect 190 875 191 876
rect 195 878 196 879
rect 274 879 280 880
rect 274 878 275 879
rect 195 876 275 878
rect 195 875 196 876
rect 190 874 196 875
rect 274 875 275 876
rect 279 875 280 879
rect 426 879 427 880
rect 431 879 432 883
rect 426 878 432 879
rect 434 879 440 880
rect 274 874 280 875
rect 338 875 344 876
rect 338 874 339 875
rect 301 872 339 874
rect 338 871 339 872
rect 343 871 344 875
rect 338 870 344 871
rect 346 875 352 876
rect 346 871 347 875
rect 351 874 352 875
rect 434 875 435 879
rect 439 878 440 879
rect 702 879 708 880
rect 702 878 703 879
rect 439 876 703 878
rect 439 875 440 876
rect 434 874 440 875
rect 702 875 703 876
rect 707 875 708 879
rect 702 874 708 875
rect 351 872 377 874
rect 351 871 352 872
rect 346 870 352 871
rect 726 871 732 872
rect 726 870 727 871
rect 612 868 727 870
rect 146 863 152 864
rect 146 862 147 863
rect 140 860 147 862
rect 140 853 142 860
rect 146 859 147 860
rect 151 862 152 863
rect 538 863 544 864
rect 612 863 614 868
rect 726 867 727 868
rect 731 867 732 871
rect 726 866 732 867
rect 538 862 539 863
rect 151 860 162 862
rect 151 859 152 860
rect 146 858 152 859
rect 160 858 162 860
rect 216 860 539 862
rect 216 858 218 860
rect 160 856 218 858
rect 338 859 344 860
rect 150 855 156 856
rect 150 851 151 855
rect 155 851 156 855
rect 150 850 156 851
rect 222 855 228 856
rect 222 851 223 855
rect 227 854 228 855
rect 230 855 236 856
rect 230 854 231 855
rect 227 852 231 854
rect 227 851 228 852
rect 222 850 228 851
rect 230 851 231 852
rect 235 851 236 855
rect 338 855 339 859
rect 343 855 344 859
rect 538 859 539 860
rect 543 859 544 863
rect 538 858 544 859
rect 338 854 344 855
rect 526 855 532 856
rect 230 850 236 851
rect 378 851 384 852
rect 166 847 172 848
rect 166 843 167 847
rect 171 843 172 847
rect 358 847 364 848
rect 358 846 359 847
rect 333 844 359 846
rect 166 842 172 843
rect 358 843 359 844
rect 363 843 364 847
rect 378 847 379 851
rect 383 847 384 851
rect 378 846 384 847
rect 386 851 392 852
rect 386 847 387 851
rect 391 850 392 851
rect 518 851 524 852
rect 518 850 519 851
rect 391 848 519 850
rect 391 847 392 848
rect 386 846 392 847
rect 518 847 519 848
rect 523 847 524 851
rect 526 851 527 855
rect 531 854 532 855
rect 624 854 626 861
rect 726 859 732 860
rect 654 855 660 856
rect 654 854 655 855
rect 531 852 626 854
rect 641 852 655 854
rect 531 851 532 852
rect 526 850 532 851
rect 654 851 655 852
rect 659 851 660 855
rect 654 850 660 851
rect 702 855 708 856
rect 702 851 703 855
rect 707 851 708 855
rect 726 855 727 859
rect 731 858 732 859
rect 766 859 772 860
rect 766 858 767 859
rect 731 856 767 858
rect 731 855 732 856
rect 726 854 732 855
rect 766 855 767 856
rect 771 855 772 859
rect 766 854 772 855
rect 702 850 708 851
rect 898 851 904 852
rect 518 846 524 847
rect 562 847 568 848
rect 358 842 364 843
rect 562 843 563 847
rect 567 846 568 847
rect 898 847 899 851
rect 903 847 904 851
rect 898 846 904 847
rect 567 844 601 846
rect 567 843 568 844
rect 562 842 568 843
rect 846 842 852 843
rect 174 840 180 841
rect 574 840 580 841
rect 174 836 175 840
rect 179 836 180 840
rect 174 835 180 836
rect 326 839 332 840
rect 326 835 327 839
rect 331 835 332 839
rect 574 836 575 840
rect 579 836 580 840
rect 326 834 332 835
rect 450 835 456 836
rect 574 835 580 836
rect 774 840 780 841
rect 774 836 775 840
rect 779 836 780 840
rect 774 835 780 836
rect 806 840 812 841
rect 806 836 807 840
rect 811 836 812 840
rect 846 838 847 842
rect 851 838 852 842
rect 846 837 852 838
rect 806 835 812 836
rect 110 833 116 834
rect 110 829 111 833
rect 115 829 116 833
rect 450 831 451 835
rect 455 831 456 835
rect 958 833 964 834
rect 450 830 456 831
rect 518 831 524 832
rect 110 828 116 829
rect 274 827 280 828
rect 274 823 275 827
rect 279 826 280 827
rect 346 827 352 828
rect 346 826 347 827
rect 279 824 347 826
rect 279 823 280 824
rect 274 822 280 823
rect 346 823 347 824
rect 351 823 352 827
rect 518 827 519 831
rect 523 827 524 831
rect 638 829 644 830
rect 518 826 524 827
rect 586 827 592 828
rect 586 826 587 827
rect 520 824 587 826
rect 346 822 352 823
rect 586 823 587 824
rect 591 823 592 827
rect 638 825 639 829
rect 643 825 644 829
rect 958 829 959 833
rect 963 829 964 833
rect 958 828 964 829
rect 638 824 644 825
rect 586 822 592 823
rect 513 820 518 822
rect 516 818 522 820
rect 594 819 600 820
rect 594 818 595 819
rect 158 816 164 817
rect 110 815 116 816
rect 110 811 111 815
rect 115 811 116 815
rect 158 812 159 816
rect 163 812 164 816
rect 158 811 164 812
rect 450 816 456 817
rect 520 816 595 818
rect 450 812 451 816
rect 455 812 456 816
rect 594 815 595 816
rect 599 815 600 819
rect 766 819 772 820
rect 594 814 600 815
rect 638 816 644 817
rect 638 812 639 816
rect 643 812 644 816
rect 766 815 767 819
rect 771 818 772 819
rect 799 819 805 820
rect 771 816 785 818
rect 771 815 772 816
rect 766 814 772 815
rect 799 815 800 819
rect 804 818 805 819
rect 804 816 817 818
rect 846 816 852 817
rect 804 815 805 816
rect 799 814 805 815
rect 846 812 847 816
rect 851 812 852 816
rect 450 811 456 812
rect 586 811 592 812
rect 110 810 116 811
rect 574 808 580 809
rect 202 807 208 808
rect 127 803 133 804
rect 127 799 128 803
rect 132 802 133 803
rect 167 803 173 804
rect 167 802 168 803
rect 132 800 168 802
rect 132 799 133 800
rect 127 798 133 799
rect 167 799 168 800
rect 172 799 173 803
rect 202 803 203 807
rect 207 806 208 807
rect 470 807 476 808
rect 207 804 254 806
rect 207 803 208 804
rect 202 802 208 803
rect 252 802 254 804
rect 382 803 388 804
rect 252 800 269 802
rect 167 798 173 799
rect 382 799 383 803
rect 387 799 388 803
rect 470 803 471 807
rect 475 803 476 807
rect 574 804 575 808
rect 579 804 580 808
rect 586 807 587 811
rect 591 807 592 811
rect 586 806 592 807
rect 630 811 636 812
rect 638 811 644 812
rect 826 811 832 812
rect 846 811 852 812
rect 958 815 964 816
rect 958 811 959 815
rect 963 811 964 815
rect 630 807 631 811
rect 635 807 636 811
rect 630 806 636 807
rect 774 808 780 809
rect 574 803 580 804
rect 774 804 775 808
rect 779 804 780 808
rect 806 808 812 809
rect 774 803 780 804
rect 470 802 476 803
rect 382 798 388 799
rect 554 799 560 800
rect 554 798 555 799
rect 416 796 555 798
rect 274 795 280 796
rect 274 791 275 795
rect 279 791 280 795
rect 274 790 280 791
rect 310 793 316 794
rect 310 789 311 793
rect 315 789 316 793
rect 416 790 418 796
rect 554 795 555 796
rect 559 795 560 799
rect 554 794 560 795
rect 738 799 744 800
rect 738 795 739 799
rect 743 798 744 799
rect 784 798 786 805
rect 806 804 807 808
rect 811 804 812 808
rect 806 803 812 804
rect 818 807 824 808
rect 818 803 819 807
rect 823 803 824 807
rect 826 807 827 811
rect 831 810 832 811
rect 958 810 964 811
rect 831 808 841 810
rect 831 807 832 808
rect 826 806 832 807
rect 818 802 824 803
rect 743 796 786 798
rect 743 795 744 796
rect 738 794 744 795
rect 834 795 840 796
rect 834 791 835 795
rect 839 791 840 795
rect 834 790 840 791
rect 854 795 860 796
rect 854 791 855 795
rect 859 794 860 795
rect 859 792 905 794
rect 859 791 860 792
rect 854 790 860 791
rect 310 788 316 789
rect 376 788 418 790
rect 488 788 566 790
rect 126 787 132 788
rect 126 783 127 787
rect 131 786 132 787
rect 167 787 173 788
rect 131 784 145 786
rect 131 783 132 784
rect 126 782 132 783
rect 167 783 168 787
rect 172 786 173 787
rect 366 787 372 788
rect 366 786 367 787
rect 172 784 181 786
rect 284 784 367 786
rect 172 783 173 784
rect 167 782 173 783
rect 284 782 286 784
rect 160 778 162 781
rect 241 780 286 782
rect 198 779 204 780
rect 198 778 199 779
rect 160 776 199 778
rect 198 775 199 776
rect 203 775 204 779
rect 198 774 204 775
rect 298 779 304 780
rect 328 779 330 784
rect 366 783 367 784
rect 371 783 372 787
rect 366 782 372 783
rect 374 787 380 788
rect 374 783 375 787
rect 379 783 380 787
rect 374 782 380 783
rect 442 787 448 788
rect 442 783 443 787
rect 447 786 448 787
rect 486 787 492 788
rect 486 786 487 787
rect 447 784 487 786
rect 447 783 448 784
rect 442 782 448 783
rect 486 783 487 784
rect 491 783 492 787
rect 564 786 566 788
rect 639 787 645 788
rect 564 784 617 786
rect 486 782 492 783
rect 626 783 632 784
rect 366 779 372 780
rect 298 775 299 779
rect 303 778 304 779
rect 366 778 367 779
rect 303 776 309 778
rect 357 776 367 778
rect 303 775 304 776
rect 298 774 304 775
rect 366 775 367 776
rect 371 775 372 779
rect 626 779 627 783
rect 631 779 632 783
rect 639 783 640 787
rect 644 786 645 787
rect 644 784 685 786
rect 848 784 850 789
rect 644 783 645 784
rect 639 782 645 783
rect 847 783 853 784
rect 626 778 632 779
rect 847 779 848 783
rect 852 779 853 783
rect 847 778 853 779
rect 366 774 372 775
rect 430 771 436 772
rect 430 767 431 771
rect 435 767 436 771
rect 511 771 517 772
rect 511 770 512 771
rect 457 769 512 770
rect 456 768 512 769
rect 430 766 436 767
rect 442 767 448 768
rect 167 763 173 764
rect 167 759 168 763
rect 172 762 173 763
rect 318 763 324 764
rect 172 760 289 762
rect 172 759 173 760
rect 318 759 319 763
rect 323 762 324 763
rect 366 763 372 764
rect 366 762 367 763
rect 323 760 367 762
rect 323 759 324 760
rect 167 758 173 759
rect 238 755 244 756
rect 238 751 239 755
rect 243 754 244 755
rect 300 754 302 759
rect 318 758 324 759
rect 366 759 367 760
rect 371 759 372 763
rect 442 763 443 767
rect 447 763 448 767
rect 442 762 448 763
rect 366 758 372 759
rect 456 758 458 768
rect 511 767 512 768
rect 516 767 517 771
rect 511 766 517 767
rect 526 771 532 772
rect 526 767 527 771
rect 531 767 532 771
rect 526 766 532 767
rect 538 771 544 772
rect 538 767 539 771
rect 543 767 544 771
rect 538 766 544 767
rect 554 771 560 772
rect 554 767 555 771
rect 559 770 560 771
rect 682 771 688 772
rect 682 770 683 771
rect 559 768 683 770
rect 559 767 560 768
rect 554 766 560 767
rect 682 767 683 768
rect 687 767 688 771
rect 682 766 688 767
rect 510 763 516 764
rect 510 759 511 763
rect 515 762 516 763
rect 626 763 632 764
rect 626 762 627 763
rect 515 760 627 762
rect 515 759 516 760
rect 510 758 516 759
rect 626 759 627 760
rect 631 759 632 763
rect 626 758 632 759
rect 818 763 824 764
rect 818 759 819 763
rect 823 762 824 763
rect 855 763 861 764
rect 855 762 856 763
rect 823 760 856 762
rect 823 759 824 760
rect 818 758 824 759
rect 855 759 856 760
rect 860 759 861 763
rect 855 758 861 759
rect 368 756 458 758
rect 828 756 850 758
rect 526 755 532 756
rect 526 754 527 755
rect 243 752 527 754
rect 243 751 244 752
rect 238 750 244 751
rect 526 751 527 752
rect 531 751 532 755
rect 526 750 532 751
rect 535 755 541 756
rect 535 751 536 755
rect 540 754 541 755
rect 550 755 556 756
rect 550 754 551 755
rect 540 752 551 754
rect 540 751 541 752
rect 535 750 541 751
rect 550 751 551 752
rect 555 754 556 755
rect 666 755 672 756
rect 666 754 667 755
rect 555 752 667 754
rect 555 751 556 752
rect 550 750 556 751
rect 666 751 667 752
rect 671 754 672 755
rect 710 755 716 756
rect 710 754 711 755
rect 671 752 711 754
rect 671 751 672 752
rect 666 750 672 751
rect 710 751 711 752
rect 715 754 716 755
rect 828 754 830 756
rect 715 752 830 754
rect 847 755 853 756
rect 715 751 716 752
rect 710 750 716 751
rect 834 751 840 752
rect 476 748 518 750
rect 358 747 364 748
rect 358 743 359 747
rect 363 746 364 747
rect 450 747 456 748
rect 450 746 451 747
rect 363 744 451 746
rect 363 743 364 744
rect 358 742 364 743
rect 450 743 451 744
rect 455 746 456 747
rect 476 747 484 748
rect 476 746 479 747
rect 455 744 479 746
rect 455 743 456 744
rect 450 742 456 743
rect 478 743 479 744
rect 483 743 484 747
rect 516 746 518 748
rect 639 747 645 748
rect 639 746 640 747
rect 516 744 640 746
rect 478 742 484 743
rect 506 743 512 744
rect 294 739 300 740
rect 294 738 295 739
rect 164 736 295 738
rect 164 729 166 736
rect 294 735 295 736
rect 299 738 300 739
rect 374 739 380 740
rect 374 738 375 739
rect 299 736 375 738
rect 299 735 300 736
rect 294 734 300 735
rect 374 735 375 736
rect 379 735 380 739
rect 506 739 507 743
rect 511 742 512 743
rect 639 743 640 744
rect 644 743 645 747
rect 639 742 645 743
rect 790 747 796 748
rect 790 743 791 747
rect 795 746 796 747
rect 822 747 828 748
rect 822 746 823 747
rect 795 744 823 746
rect 795 743 796 744
rect 790 742 796 743
rect 822 743 823 744
rect 827 743 828 747
rect 834 747 835 751
rect 839 747 840 751
rect 847 751 848 755
rect 852 751 853 755
rect 847 750 853 751
rect 834 746 840 747
rect 848 745 850 750
rect 855 747 864 748
rect 822 742 828 743
rect 855 743 856 747
rect 863 743 864 747
rect 855 742 864 743
rect 866 747 872 748
rect 866 743 867 747
rect 871 743 872 747
rect 866 742 872 743
rect 926 747 932 748
rect 926 743 927 747
rect 931 743 932 747
rect 926 742 932 743
rect 511 740 598 742
rect 511 739 512 740
rect 506 738 512 739
rect 594 739 600 740
rect 516 736 529 738
rect 545 736 554 738
rect 374 734 380 735
rect 514 735 520 736
rect 198 731 204 732
rect 198 730 199 731
rect 177 728 199 730
rect 198 727 199 728
rect 203 727 204 731
rect 198 726 204 727
rect 230 731 236 732
rect 230 727 231 731
rect 235 727 236 731
rect 514 731 515 735
rect 519 731 520 735
rect 514 730 520 731
rect 550 735 556 736
rect 550 731 551 735
rect 555 731 556 735
rect 550 730 556 731
rect 562 735 568 736
rect 562 731 563 735
rect 567 731 568 735
rect 594 735 595 739
rect 599 735 600 739
rect 594 734 600 735
rect 682 739 688 740
rect 682 735 683 739
rect 687 738 688 739
rect 799 739 805 740
rect 799 738 800 739
rect 687 736 800 738
rect 687 735 688 736
rect 682 734 688 735
rect 799 735 800 736
rect 804 735 805 739
rect 799 734 805 735
rect 562 730 568 731
rect 684 729 686 734
rect 710 731 716 732
rect 710 730 711 731
rect 697 728 711 730
rect 230 726 236 727
rect 710 727 711 728
rect 715 727 716 731
rect 766 731 772 732
rect 766 730 767 731
rect 757 728 767 730
rect 710 726 716 727
rect 766 727 767 728
rect 771 727 772 731
rect 766 726 772 727
rect 488 724 518 726
rect 314 723 320 724
rect 314 719 315 723
rect 319 719 320 723
rect 374 719 380 720
rect 314 718 320 719
rect 350 718 356 719
rect 374 718 375 719
rect 134 716 140 717
rect 134 712 135 716
rect 139 712 140 716
rect 278 716 284 717
rect 302 716 308 717
rect 149 712 169 714
rect 278 712 279 716
rect 283 712 284 716
rect 134 711 140 712
rect 278 711 284 712
rect 290 715 296 716
rect 290 711 291 715
rect 295 711 296 715
rect 302 712 303 716
rect 307 712 308 716
rect 316 713 318 718
rect 326 716 332 717
rect 302 711 308 712
rect 326 712 327 716
rect 331 712 332 716
rect 326 711 332 712
rect 338 715 344 716
rect 338 711 339 715
rect 343 711 344 715
rect 350 714 351 718
rect 355 714 356 718
rect 365 716 375 718
rect 374 715 375 716
rect 379 715 380 719
rect 414 718 420 719
rect 374 714 380 715
rect 382 716 388 717
rect 350 713 356 714
rect 382 712 383 716
rect 387 712 388 716
rect 406 715 412 716
rect 406 714 407 715
rect 397 712 407 714
rect 382 711 388 712
rect 406 711 407 712
rect 411 711 412 715
rect 414 714 415 718
rect 419 714 420 718
rect 414 713 420 714
rect 438 716 444 717
rect 462 716 468 717
rect 290 710 296 711
rect 338 710 344 711
rect 406 710 412 711
rect 424 710 426 713
rect 438 712 439 716
rect 443 712 444 716
rect 438 711 444 712
rect 450 715 456 716
rect 450 711 451 715
rect 455 711 456 715
rect 462 712 463 716
rect 467 712 468 716
rect 488 714 490 724
rect 506 719 512 720
rect 477 712 490 714
rect 494 718 500 719
rect 494 714 495 718
rect 499 714 500 718
rect 506 715 507 719
rect 511 715 512 719
rect 506 714 512 715
rect 516 714 518 724
rect 918 723 924 724
rect 918 719 919 723
rect 923 722 924 723
rect 1011 723 1017 724
rect 1011 722 1012 723
rect 923 720 1012 722
rect 923 719 924 720
rect 918 718 924 719
rect 1011 719 1012 720
rect 1016 719 1017 723
rect 1011 718 1017 719
rect 654 716 660 717
rect 494 713 500 714
rect 516 712 537 714
rect 654 712 655 716
rect 659 712 660 716
rect 798 716 804 717
rect 669 712 689 714
rect 798 712 799 716
rect 803 712 804 716
rect 823 715 829 716
rect 823 714 824 715
rect 813 712 824 714
rect 462 711 468 712
rect 654 711 660 712
rect 798 711 804 712
rect 823 711 824 712
rect 828 714 829 715
rect 834 715 840 716
rect 834 714 835 715
rect 828 712 835 714
rect 828 711 829 712
rect 450 710 456 711
rect 823 710 829 711
rect 834 711 835 712
rect 839 711 840 715
rect 834 710 840 711
rect 110 709 116 710
rect 110 705 111 709
rect 115 705 116 709
rect 110 704 116 705
rect 174 708 180 709
rect 424 708 434 710
rect 958 709 964 710
rect 542 708 548 709
rect 174 704 175 708
rect 179 704 180 708
rect 142 703 148 704
rect 174 703 180 704
rect 286 703 292 704
rect 142 699 143 703
rect 147 699 148 703
rect 142 698 148 699
rect 286 699 287 703
rect 291 699 292 703
rect 358 703 364 704
rect 286 698 292 699
rect 263 695 269 696
rect 110 691 116 692
rect 110 687 111 691
rect 115 687 116 691
rect 263 691 264 695
rect 268 694 269 695
rect 312 694 314 701
rect 268 692 314 694
rect 336 694 338 701
rect 358 699 359 703
rect 363 699 364 703
rect 358 698 364 699
rect 390 703 396 704
rect 390 699 391 703
rect 395 699 396 703
rect 390 698 396 699
rect 422 703 428 704
rect 422 699 423 703
rect 427 699 428 703
rect 432 702 434 708
rect 486 707 492 708
rect 446 703 452 704
rect 446 702 447 703
rect 432 700 447 702
rect 422 698 428 699
rect 446 699 447 700
rect 451 699 452 703
rect 486 703 487 707
rect 491 706 492 707
rect 491 704 505 706
rect 542 704 543 708
rect 547 704 548 708
rect 694 708 700 709
rect 694 704 695 708
rect 699 704 700 708
rect 846 708 852 709
rect 846 704 847 708
rect 851 704 852 708
rect 958 705 959 709
rect 963 705 964 709
rect 958 704 964 705
rect 491 703 492 704
rect 542 703 548 704
rect 662 703 668 704
rect 694 703 700 704
rect 806 703 812 704
rect 846 703 852 704
rect 486 702 492 703
rect 446 698 452 699
rect 472 698 474 701
rect 486 699 492 700
rect 486 698 487 699
rect 472 696 487 698
rect 406 695 412 696
rect 406 694 407 695
rect 336 692 407 694
rect 268 691 269 692
rect 263 690 269 691
rect 406 691 407 692
rect 411 691 412 695
rect 486 695 487 696
rect 491 695 492 699
rect 662 699 663 703
rect 667 699 668 703
rect 662 698 668 699
rect 806 699 807 703
rect 811 699 812 703
rect 806 698 812 699
rect 486 694 492 695
rect 542 694 548 695
rect 406 690 412 691
rect 542 690 543 694
rect 547 690 548 694
rect 542 689 548 690
rect 846 691 852 692
rect 110 686 116 687
rect 846 687 847 691
rect 851 687 852 691
rect 846 686 852 687
rect 958 691 964 692
rect 958 687 959 691
rect 963 687 964 691
rect 958 686 964 687
rect 134 684 140 685
rect 134 680 135 684
rect 139 680 140 684
rect 278 684 284 685
rect 134 679 140 680
rect 174 682 180 683
rect 174 678 175 682
rect 179 678 180 682
rect 278 680 279 684
rect 283 680 284 684
rect 278 679 284 680
rect 302 684 308 685
rect 302 680 303 684
rect 307 680 308 684
rect 302 679 308 680
rect 326 684 332 685
rect 326 680 327 684
rect 331 680 332 684
rect 326 679 332 680
rect 350 684 356 685
rect 350 680 351 684
rect 355 680 356 684
rect 350 679 356 680
rect 382 684 388 685
rect 382 680 383 684
rect 387 680 388 684
rect 382 679 388 680
rect 414 684 420 685
rect 414 680 415 684
rect 419 680 420 684
rect 414 679 420 680
rect 438 684 444 685
rect 438 680 439 684
rect 443 680 444 684
rect 438 679 444 680
rect 462 684 468 685
rect 462 680 463 684
rect 467 680 468 684
rect 462 679 468 680
rect 494 684 500 685
rect 494 680 495 684
rect 499 680 500 684
rect 494 679 500 680
rect 654 684 660 685
rect 654 680 655 684
rect 659 680 660 684
rect 798 684 804 685
rect 654 679 660 680
rect 694 682 700 683
rect 174 677 180 678
rect 694 678 695 682
rect 699 678 700 682
rect 798 680 799 684
rect 803 680 804 684
rect 798 679 804 680
rect 938 679 944 680
rect 938 678 939 679
rect 694 677 700 678
rect 808 676 841 678
rect 880 676 939 678
rect 150 675 156 676
rect 150 671 151 675
rect 155 674 156 675
rect 358 675 364 676
rect 358 674 359 675
rect 155 673 229 674
rect 233 673 359 674
rect 155 672 230 673
rect 155 671 156 672
rect 150 670 156 671
rect 228 670 230 672
rect 232 672 359 673
rect 232 670 234 672
rect 358 671 359 672
rect 363 674 364 675
rect 562 675 568 676
rect 562 674 563 675
rect 363 672 563 674
rect 363 671 364 672
rect 358 670 364 671
rect 562 671 563 672
rect 567 674 568 675
rect 758 675 764 676
rect 567 672 749 674
rect 567 671 568 672
rect 562 670 568 671
rect 758 671 759 675
rect 763 674 764 675
rect 808 674 810 676
rect 763 672 810 674
rect 763 671 764 672
rect 758 670 764 671
rect 834 671 840 672
rect 228 668 234 670
rect 142 667 148 668
rect 142 663 143 667
rect 147 666 148 667
rect 318 667 324 668
rect 318 666 319 667
rect 147 664 319 666
rect 147 663 148 664
rect 142 662 148 663
rect 318 663 319 664
rect 323 666 324 667
rect 327 667 333 668
rect 327 666 328 667
rect 323 664 328 666
rect 323 663 324 664
rect 318 662 324 663
rect 327 663 328 664
rect 332 663 333 667
rect 327 662 333 663
rect 471 667 477 668
rect 471 663 472 667
rect 476 666 477 667
rect 670 667 676 668
rect 670 666 671 667
rect 476 664 671 666
rect 476 663 477 664
rect 471 662 477 663
rect 670 663 671 664
rect 675 663 676 667
rect 834 667 835 671
rect 839 670 840 671
rect 880 670 882 676
rect 938 675 939 676
rect 943 675 944 679
rect 938 674 944 675
rect 839 668 882 670
rect 839 667 840 668
rect 834 666 840 667
rect 670 662 676 663
rect 806 663 812 664
rect 662 659 668 660
rect 662 658 663 659
rect 616 656 663 658
rect 294 651 300 652
rect 294 650 295 651
rect 264 648 295 650
rect 264 646 266 648
rect 294 647 295 648
rect 299 650 300 651
rect 594 651 600 652
rect 299 648 470 650
rect 299 647 300 648
rect 294 646 300 647
rect 466 647 472 648
rect 144 644 266 646
rect 144 641 146 644
rect 264 641 266 644
rect 274 643 280 644
rect 255 639 261 640
rect 255 638 256 639
rect 225 636 256 638
rect 255 635 256 636
rect 260 635 261 639
rect 274 639 275 643
rect 279 639 280 643
rect 274 638 280 639
rect 327 643 333 644
rect 327 639 328 643
rect 332 642 333 643
rect 466 643 467 647
rect 471 643 472 647
rect 594 647 595 651
rect 599 650 600 651
rect 616 650 618 656
rect 662 655 663 656
rect 667 655 668 659
rect 806 659 807 663
rect 811 662 812 663
rect 818 663 824 664
rect 818 662 819 663
rect 811 660 819 662
rect 811 659 812 660
rect 806 658 812 659
rect 818 659 819 660
rect 823 662 824 663
rect 912 662 914 669
rect 823 660 914 662
rect 823 659 824 660
rect 818 658 824 659
rect 662 654 668 655
rect 638 651 644 652
rect 599 648 621 650
rect 599 647 600 648
rect 594 646 600 647
rect 466 642 472 643
rect 618 643 624 644
rect 332 640 349 642
rect 332 639 333 640
rect 327 638 333 639
rect 566 639 572 640
rect 566 638 567 639
rect 509 636 567 638
rect 255 634 261 635
rect 334 635 340 636
rect 334 634 335 635
rect 317 632 335 634
rect 262 631 268 632
rect 262 630 263 631
rect 165 628 263 630
rect 262 627 263 628
rect 267 627 268 631
rect 334 631 335 632
rect 339 631 340 635
rect 334 630 340 631
rect 430 635 436 636
rect 430 631 431 635
rect 435 634 436 635
rect 471 635 477 636
rect 471 634 472 635
rect 435 632 472 634
rect 435 631 436 632
rect 430 630 436 631
rect 471 631 472 632
rect 476 631 477 635
rect 566 635 567 636
rect 571 635 572 639
rect 618 639 619 643
rect 623 642 624 643
rect 632 642 634 649
rect 638 647 639 651
rect 643 650 644 651
rect 830 651 836 652
rect 830 650 831 651
rect 643 648 714 650
rect 643 647 644 648
rect 638 646 644 647
rect 678 643 684 644
rect 678 642 679 643
rect 623 640 634 642
rect 649 640 679 642
rect 623 639 624 640
rect 618 638 624 639
rect 678 639 679 640
rect 683 639 684 643
rect 712 641 714 648
rect 804 648 831 650
rect 804 641 806 648
rect 830 647 831 648
rect 835 647 836 651
rect 830 646 836 647
rect 810 643 816 644
rect 678 638 684 639
rect 810 639 811 643
rect 815 639 816 643
rect 810 638 816 639
rect 823 643 829 644
rect 823 639 824 643
rect 828 642 829 643
rect 828 640 885 642
rect 828 639 829 640
rect 823 638 829 639
rect 566 634 572 635
rect 606 635 612 636
rect 471 630 477 631
rect 606 631 607 635
rect 611 631 612 635
rect 606 630 612 631
rect 798 631 804 632
rect 262 626 268 627
rect 302 628 308 629
rect 558 628 564 629
rect 302 624 303 628
rect 307 624 308 628
rect 302 623 308 624
rect 454 627 460 628
rect 454 623 455 627
rect 459 623 460 627
rect 558 624 559 628
rect 563 624 564 628
rect 558 623 564 624
rect 582 628 588 629
rect 582 624 583 628
rect 587 624 588 628
rect 582 623 588 624
rect 774 628 780 629
rect 774 624 775 628
rect 779 624 780 628
rect 798 627 799 631
rect 803 630 804 631
rect 803 628 817 630
rect 838 628 844 629
rect 803 627 804 628
rect 798 626 804 627
rect 774 623 780 624
rect 838 624 839 628
rect 843 624 844 628
rect 838 623 844 624
rect 926 628 932 629
rect 926 624 927 628
rect 931 624 932 628
rect 926 623 932 624
rect 454 622 460 623
rect 110 621 116 622
rect 110 617 111 621
rect 115 617 116 621
rect 110 616 116 617
rect 158 621 164 622
rect 158 617 159 621
rect 163 617 164 621
rect 958 621 964 622
rect 158 616 164 617
rect 646 617 652 618
rect 510 615 516 616
rect 510 614 511 615
rect 360 612 511 614
rect 230 611 236 612
rect 230 607 231 611
rect 235 610 236 611
rect 274 611 280 612
rect 274 610 275 611
rect 235 608 275 610
rect 235 607 236 608
rect 230 606 236 607
rect 274 607 275 608
rect 279 607 280 611
rect 274 606 280 607
rect 358 611 364 612
rect 358 607 359 611
rect 363 607 364 611
rect 510 611 511 612
rect 515 611 516 615
rect 510 610 516 611
rect 538 615 544 616
rect 538 611 539 615
rect 543 614 544 615
rect 543 612 578 614
rect 646 613 647 617
rect 651 613 652 617
rect 958 617 959 621
rect 963 617 964 621
rect 958 616 964 617
rect 646 612 652 613
rect 543 611 544 612
rect 538 610 544 611
rect 358 606 364 607
rect 550 607 556 608
rect 158 604 164 605
rect 110 603 116 604
rect 110 599 111 603
rect 115 599 116 603
rect 158 600 159 604
rect 163 600 164 604
rect 158 599 164 600
rect 286 604 292 605
rect 286 600 287 604
rect 291 600 292 604
rect 550 603 551 607
rect 555 606 556 607
rect 566 607 572 608
rect 566 606 567 607
rect 555 604 567 606
rect 555 603 556 604
rect 550 602 556 603
rect 566 603 567 604
rect 571 603 572 607
rect 576 606 578 612
rect 638 607 644 608
rect 638 606 639 607
rect 576 604 639 606
rect 566 602 572 603
rect 638 603 639 604
rect 643 603 644 607
rect 782 607 788 608
rect 638 602 644 603
rect 646 604 652 605
rect 646 600 647 604
rect 651 600 652 604
rect 782 603 783 607
rect 787 603 788 607
rect 782 602 788 603
rect 822 604 828 605
rect 286 599 292 600
rect 478 599 484 600
rect 646 599 652 600
rect 822 600 823 604
rect 827 600 828 604
rect 880 604 937 606
rect 822 599 828 600
rect 866 599 872 600
rect 110 598 116 599
rect 326 595 332 596
rect 198 591 204 592
rect 167 587 173 588
rect 167 583 168 587
rect 172 586 173 587
rect 198 587 199 591
rect 203 590 204 591
rect 278 591 284 592
rect 278 590 279 591
rect 203 588 279 590
rect 203 587 204 588
rect 198 586 204 587
rect 278 587 279 588
rect 283 587 284 591
rect 326 591 327 595
rect 331 594 332 595
rect 478 595 479 599
rect 483 595 484 599
rect 478 594 484 595
rect 558 596 564 597
rect 582 596 588 597
rect 774 596 780 597
rect 331 592 382 594
rect 331 591 332 592
rect 326 590 332 591
rect 380 590 382 592
rect 558 592 559 596
rect 563 592 564 596
rect 558 591 564 592
rect 570 595 576 596
rect 570 591 571 595
rect 575 591 576 595
rect 582 592 583 596
rect 587 592 588 596
rect 582 591 588 592
rect 594 595 600 596
rect 594 591 595 595
rect 599 591 600 595
rect 570 590 576 591
rect 594 590 600 591
rect 604 592 633 594
rect 774 592 775 596
rect 779 592 780 596
rect 798 595 804 596
rect 798 594 799 595
rect 789 592 799 594
rect 380 588 397 590
rect 278 586 284 587
rect 551 587 557 588
rect 172 584 202 586
rect 172 583 173 584
rect 167 582 173 583
rect 382 583 388 584
rect 382 579 383 583
rect 387 582 388 583
rect 551 583 552 587
rect 556 586 557 587
rect 604 586 606 592
rect 774 591 780 592
rect 798 591 799 592
rect 803 591 804 595
rect 866 595 867 599
rect 871 598 872 599
rect 880 598 882 604
rect 958 603 964 604
rect 958 599 959 603
rect 963 599 964 603
rect 958 598 964 599
rect 871 596 882 598
rect 926 596 932 597
rect 871 595 872 596
rect 866 594 872 595
rect 926 592 927 596
rect 931 592 932 596
rect 926 591 932 592
rect 938 595 944 596
rect 938 591 939 595
rect 943 591 944 595
rect 798 590 804 591
rect 938 590 944 591
rect 556 584 606 586
rect 790 587 797 588
rect 556 583 557 584
rect 551 582 557 583
rect 790 583 791 587
rect 796 583 797 587
rect 790 582 797 583
rect 387 580 405 582
rect 438 581 444 582
rect 387 579 388 580
rect 382 578 388 579
rect 438 577 439 581
rect 443 577 444 581
rect 438 576 444 577
rect 294 575 301 576
rect 255 571 261 572
rect 167 567 173 568
rect 167 566 168 567
rect 161 564 168 566
rect 134 563 140 564
rect 134 559 135 563
rect 139 559 140 563
rect 134 558 140 559
rect 146 563 152 564
rect 146 559 147 563
rect 151 559 152 563
rect 167 563 168 564
rect 172 563 173 567
rect 255 567 256 571
rect 260 570 261 571
rect 278 571 284 572
rect 260 569 273 570
rect 260 568 274 569
rect 260 567 261 568
rect 255 566 261 567
rect 167 562 173 563
rect 146 558 152 559
rect 184 554 186 565
rect 238 563 244 564
rect 238 559 239 563
rect 243 559 244 563
rect 272 562 274 568
rect 278 567 279 571
rect 283 570 284 571
rect 294 571 295 575
rect 300 574 301 575
rect 350 575 356 576
rect 300 572 309 574
rect 300 571 301 572
rect 294 570 301 571
rect 350 571 351 575
rect 355 574 356 575
rect 519 575 525 576
rect 355 572 446 574
rect 355 571 356 572
rect 350 570 356 571
rect 283 569 289 570
rect 283 568 290 569
rect 283 567 284 568
rect 278 566 284 567
rect 288 566 290 568
rect 376 568 395 570
rect 376 566 378 568
rect 288 564 378 566
rect 391 567 397 568
rect 382 563 388 564
rect 382 562 383 563
rect 272 560 383 562
rect 238 558 244 559
rect 382 559 383 560
rect 387 559 388 563
rect 391 563 392 567
rect 396 563 397 567
rect 391 562 397 563
rect 410 567 416 568
rect 410 563 411 567
rect 415 566 416 567
rect 444 566 446 572
rect 519 571 520 575
rect 524 574 525 575
rect 670 575 676 576
rect 524 572 625 574
rect 524 571 525 572
rect 519 570 525 571
rect 670 571 671 575
rect 675 574 676 575
rect 794 575 800 576
rect 675 572 693 574
rect 675 571 676 572
rect 670 570 676 571
rect 794 571 795 575
rect 799 574 800 575
rect 814 575 820 576
rect 814 574 815 575
rect 799 572 815 574
rect 799 571 800 572
rect 794 570 800 571
rect 814 571 815 572
rect 819 571 820 575
rect 846 575 852 576
rect 814 570 820 571
rect 830 571 836 572
rect 830 570 831 571
rect 454 567 460 568
rect 454 566 455 567
rect 415 564 437 566
rect 444 564 455 566
rect 415 563 416 564
rect 410 562 416 563
rect 454 563 455 564
rect 459 563 460 567
rect 495 567 501 568
rect 495 566 496 567
rect 485 564 496 566
rect 454 562 460 563
rect 495 563 496 564
rect 500 563 501 567
rect 640 566 642 569
rect 825 568 831 570
rect 830 567 831 568
rect 835 567 836 571
rect 846 571 847 575
rect 851 574 852 575
rect 866 575 872 576
rect 866 574 867 575
rect 851 572 867 574
rect 851 571 852 572
rect 846 570 852 571
rect 866 571 867 572
rect 871 571 872 575
rect 866 570 872 571
rect 878 571 884 572
rect 830 566 836 567
rect 878 567 879 571
rect 883 570 884 571
rect 883 568 905 570
rect 883 567 884 568
rect 878 566 884 567
rect 636 564 642 566
rect 495 562 501 563
rect 550 563 556 564
rect 382 558 388 559
rect 482 559 488 560
rect 295 555 301 556
rect 295 554 296 555
rect 184 552 296 554
rect 295 551 296 552
rect 300 554 301 555
rect 482 555 483 559
rect 487 555 488 559
rect 550 559 551 563
rect 555 562 556 563
rect 636 562 638 564
rect 555 560 638 562
rect 810 563 816 564
rect 555 559 556 560
rect 550 558 556 559
rect 810 559 811 563
rect 815 562 816 563
rect 946 563 952 564
rect 946 562 947 563
rect 815 560 947 562
rect 815 559 816 560
rect 810 558 816 559
rect 946 559 947 560
rect 951 559 952 563
rect 946 558 952 559
rect 482 554 488 555
rect 570 555 576 556
rect 300 552 321 554
rect 300 551 301 552
rect 295 550 301 551
rect 319 546 321 552
rect 454 551 460 552
rect 416 546 418 549
rect 454 547 455 551
rect 459 550 460 551
rect 570 551 571 555
rect 575 551 576 555
rect 570 550 576 551
rect 710 555 716 556
rect 710 551 711 555
rect 715 554 716 555
rect 830 555 836 556
rect 830 554 831 555
rect 715 552 831 554
rect 715 551 716 552
rect 710 550 716 551
rect 830 551 831 552
rect 835 554 836 555
rect 870 555 876 556
rect 870 554 871 555
rect 835 552 871 554
rect 835 551 836 552
rect 830 550 836 551
rect 870 551 871 552
rect 875 551 876 555
rect 870 550 876 551
rect 459 548 574 550
rect 459 547 460 548
rect 319 544 418 546
rect 238 543 244 544
rect 238 539 239 543
rect 243 542 244 543
rect 428 542 430 547
rect 454 546 460 547
rect 846 547 852 548
rect 846 546 847 547
rect 808 544 847 546
rect 791 543 797 544
rect 243 540 370 542
rect 428 540 454 542
rect 243 539 244 540
rect 238 538 244 539
rect 368 539 376 540
rect 368 538 371 539
rect 79 535 85 536
rect 79 531 80 535
rect 84 534 85 535
rect 167 535 173 536
rect 167 534 168 535
rect 84 532 168 534
rect 84 531 85 532
rect 79 530 85 531
rect 167 531 168 532
rect 172 531 173 535
rect 167 530 173 531
rect 358 535 364 536
rect 358 531 359 535
rect 363 531 364 535
rect 370 535 371 538
rect 375 535 376 539
rect 370 534 376 535
rect 390 539 396 540
rect 390 535 391 539
rect 395 538 396 539
rect 428 538 430 540
rect 395 536 430 538
rect 452 538 454 540
rect 614 539 620 540
rect 614 538 615 539
rect 452 536 615 538
rect 395 535 396 536
rect 390 534 396 535
rect 452 533 454 536
rect 614 535 615 536
rect 619 535 620 539
rect 791 539 792 543
rect 796 542 797 543
rect 796 540 802 542
rect 808 541 810 544
rect 846 543 847 544
rect 851 543 852 547
rect 846 542 852 543
rect 796 539 797 540
rect 791 538 797 539
rect 614 534 620 535
rect 358 530 364 531
rect 391 531 397 532
rect 391 530 392 531
rect 385 528 392 530
rect 391 527 392 528
rect 396 530 397 531
rect 438 531 444 532
rect 438 530 439 531
rect 396 528 439 530
rect 396 527 397 528
rect 391 526 397 527
rect 438 527 439 528
rect 443 527 444 531
rect 438 526 444 527
rect 466 531 472 532
rect 466 527 467 531
rect 471 527 472 531
rect 466 526 472 527
rect 482 531 488 532
rect 482 527 483 531
rect 487 527 488 531
rect 800 530 802 540
rect 838 539 844 540
rect 838 538 839 539
rect 821 536 839 538
rect 838 535 839 536
rect 843 535 844 539
rect 838 534 844 535
rect 906 531 912 532
rect 906 530 907 531
rect 800 528 907 530
rect 482 526 488 527
rect 490 527 496 528
rect 490 523 491 527
rect 495 526 496 527
rect 782 527 788 528
rect 495 524 630 526
rect 495 523 496 524
rect 490 522 496 523
rect 142 519 148 520
rect 142 515 143 519
rect 147 518 148 519
rect 550 519 556 520
rect 147 516 210 518
rect 147 515 148 516
rect 142 514 148 515
rect 138 511 144 512
rect 138 507 139 511
rect 143 507 144 511
rect 167 511 173 512
rect 167 510 168 511
rect 153 508 168 510
rect 138 506 144 507
rect 167 507 168 508
rect 172 507 173 511
rect 208 509 210 516
rect 550 515 551 519
rect 555 518 556 519
rect 582 519 588 520
rect 582 518 583 519
rect 555 516 561 518
rect 577 516 583 518
rect 555 515 556 516
rect 550 514 556 515
rect 582 515 583 516
rect 587 515 588 519
rect 606 519 612 520
rect 606 518 607 519
rect 597 516 607 518
rect 582 514 588 515
rect 606 515 607 516
rect 611 515 612 519
rect 628 517 630 524
rect 762 523 768 524
rect 762 519 763 523
rect 767 522 768 523
rect 782 523 783 527
rect 787 523 788 527
rect 906 527 907 528
rect 911 527 912 531
rect 906 526 912 527
rect 782 522 788 523
rect 870 523 876 524
rect 767 520 829 522
rect 767 519 768 520
rect 762 518 768 519
rect 606 514 612 515
rect 848 514 850 521
rect 870 519 871 523
rect 875 519 876 523
rect 870 518 876 519
rect 878 515 884 516
rect 878 514 879 515
rect 848 512 879 514
rect 370 511 376 512
rect 167 506 173 507
rect 370 507 371 511
rect 375 510 376 511
rect 422 511 428 512
rect 422 510 423 511
rect 375 508 423 510
rect 375 507 376 508
rect 370 506 376 507
rect 422 507 423 508
rect 427 510 428 511
rect 519 511 525 512
rect 519 510 520 511
rect 427 508 520 510
rect 427 507 428 508
rect 422 506 428 507
rect 519 507 520 508
rect 524 507 525 511
rect 519 506 525 507
rect 794 511 800 512
rect 794 507 795 511
rect 799 507 800 511
rect 830 511 836 512
rect 794 506 800 507
rect 810 507 816 508
rect 310 503 316 504
rect 310 499 311 503
rect 315 499 316 503
rect 310 498 316 499
rect 686 503 692 504
rect 686 499 687 503
rect 691 502 692 503
rect 710 503 716 504
rect 710 502 711 503
rect 691 500 711 502
rect 691 499 692 500
rect 686 498 692 499
rect 710 499 711 500
rect 715 499 716 503
rect 810 503 811 507
rect 815 503 816 507
rect 830 507 831 511
rect 835 507 836 511
rect 878 511 879 512
rect 883 511 884 515
rect 878 510 884 511
rect 830 506 836 507
rect 810 502 816 503
rect 789 500 814 502
rect 710 498 716 499
rect 870 499 876 500
rect 254 496 260 497
rect 278 496 284 497
rect 302 496 308 497
rect 174 495 180 496
rect 174 491 175 495
rect 179 491 180 495
rect 254 492 255 496
rect 259 492 260 496
rect 254 491 260 492
rect 266 495 272 496
rect 266 491 267 495
rect 271 491 272 495
rect 278 492 279 496
rect 283 492 284 496
rect 278 491 284 492
rect 290 495 296 496
rect 290 491 291 495
rect 295 491 296 495
rect 302 492 303 496
rect 307 492 308 496
rect 312 493 314 498
rect 326 496 332 497
rect 302 491 308 492
rect 326 492 327 496
rect 331 492 332 496
rect 340 496 373 498
rect 518 496 524 497
rect 702 496 708 497
rect 340 493 342 496
rect 326 491 332 492
rect 518 492 519 496
rect 523 492 524 496
rect 551 495 557 496
rect 551 494 552 495
rect 533 492 552 494
rect 518 491 524 492
rect 551 491 552 492
rect 556 491 557 495
rect 174 490 180 491
rect 266 490 272 491
rect 290 490 296 491
rect 551 490 557 491
rect 626 495 632 496
rect 626 491 627 495
rect 631 491 632 495
rect 702 492 703 496
rect 707 492 708 496
rect 712 493 714 498
rect 750 496 756 497
rect 702 491 708 492
rect 750 492 751 496
rect 755 492 756 496
rect 750 491 756 492
rect 762 495 768 496
rect 762 491 763 495
rect 767 491 768 495
rect 870 495 871 499
rect 875 495 876 499
rect 870 494 876 495
rect 626 490 632 491
rect 762 490 768 491
rect 110 489 116 490
rect 958 489 964 490
rect 110 485 111 489
rect 115 485 116 489
rect 110 484 116 485
rect 150 488 156 489
rect 378 488 384 489
rect 574 488 580 489
rect 150 484 151 488
rect 155 484 156 488
rect 318 487 324 488
rect 318 486 319 487
rect 313 484 319 486
rect 150 483 156 484
rect 278 483 284 484
rect 278 482 279 483
rect 265 480 279 482
rect 278 479 279 480
rect 283 479 284 483
rect 302 483 308 484
rect 302 482 303 483
rect 289 480 303 482
rect 278 478 284 479
rect 302 479 303 480
rect 307 479 308 483
rect 318 483 319 484
rect 323 483 324 487
rect 350 487 356 488
rect 350 486 351 487
rect 337 484 351 486
rect 318 482 324 483
rect 350 483 351 484
rect 355 483 356 487
rect 378 484 379 488
rect 383 484 384 488
rect 378 483 384 484
rect 430 487 436 488
rect 430 483 431 487
rect 435 486 436 487
rect 458 487 464 488
rect 458 486 459 487
rect 435 484 459 486
rect 435 483 436 484
rect 350 482 356 483
rect 430 482 436 483
rect 458 483 459 484
rect 463 483 464 487
rect 458 482 464 483
rect 466 487 472 488
rect 466 483 467 487
rect 471 486 472 487
rect 471 484 529 486
rect 574 484 575 488
rect 579 484 580 488
rect 471 483 472 484
rect 574 483 580 484
rect 678 487 684 488
rect 678 483 679 487
rect 683 486 684 487
rect 683 484 713 486
rect 958 485 959 489
rect 963 485 964 489
rect 958 484 964 485
rect 683 483 684 484
rect 466 482 472 483
rect 678 482 684 483
rect 302 478 308 479
rect 446 479 452 480
rect 446 478 447 479
rect 441 476 447 478
rect 446 475 447 476
rect 451 478 452 479
rect 490 479 496 480
rect 490 478 491 479
rect 451 476 491 478
rect 451 475 452 476
rect 446 474 452 475
rect 490 475 491 476
rect 495 475 496 479
rect 490 474 496 475
rect 574 474 580 475
rect 110 471 116 472
rect 110 467 111 471
rect 115 467 116 471
rect 574 470 575 474
rect 579 470 580 474
rect 760 474 762 481
rect 910 479 916 480
rect 910 478 911 479
rect 792 476 911 478
rect 782 475 788 476
rect 782 474 783 475
rect 760 472 783 474
rect 782 471 783 472
rect 787 471 788 475
rect 782 470 788 471
rect 110 466 116 467
rect 378 469 384 470
rect 574 469 580 470
rect 378 465 379 469
rect 383 465 384 469
rect 774 467 780 468
rect 254 464 260 465
rect 150 462 156 463
rect 150 458 151 462
rect 155 458 156 462
rect 254 460 255 464
rect 259 460 260 464
rect 254 459 260 460
rect 278 464 284 465
rect 278 460 279 464
rect 283 460 284 464
rect 278 459 284 460
rect 302 464 308 465
rect 302 460 303 464
rect 307 460 308 464
rect 302 459 308 460
rect 326 464 332 465
rect 378 464 384 465
rect 518 464 524 465
rect 326 460 327 464
rect 331 460 332 464
rect 326 459 332 460
rect 518 460 519 464
rect 523 460 524 464
rect 518 459 524 460
rect 702 464 708 465
rect 702 460 703 464
rect 707 460 708 464
rect 702 459 708 460
rect 750 464 756 465
rect 750 460 751 464
rect 755 460 756 464
rect 774 463 775 467
rect 779 466 780 467
rect 792 466 794 476
rect 910 475 911 476
rect 915 475 916 479
rect 910 474 916 475
rect 958 471 964 472
rect 958 467 959 471
rect 963 467 964 471
rect 958 466 964 467
rect 779 464 794 466
rect 846 465 852 466
rect 779 463 780 464
rect 774 462 780 463
rect 846 461 847 465
rect 851 461 852 465
rect 846 460 852 461
rect 750 459 756 460
rect 762 459 768 460
rect 150 457 156 458
rect 438 455 444 456
rect 151 451 157 452
rect 151 447 152 451
rect 156 450 157 451
rect 204 450 206 453
rect 230 451 236 452
rect 230 450 231 451
rect 156 448 231 450
rect 156 447 157 448
rect 151 446 157 447
rect 230 447 231 448
rect 235 447 236 451
rect 438 451 439 455
rect 443 454 444 455
rect 495 455 501 456
rect 495 454 496 455
rect 443 452 496 454
rect 443 451 444 452
rect 438 450 444 451
rect 495 451 496 452
rect 500 454 501 455
rect 582 455 588 456
rect 582 454 583 455
rect 500 452 583 454
rect 500 451 501 452
rect 495 450 501 451
rect 582 451 583 452
rect 587 451 588 455
rect 762 455 763 459
rect 767 458 768 459
rect 834 459 840 460
rect 834 458 835 459
rect 767 456 835 458
rect 767 455 768 456
rect 762 454 768 455
rect 834 455 835 456
rect 839 458 840 459
rect 839 456 853 458
rect 839 455 840 456
rect 834 454 840 455
rect 910 455 916 456
rect 910 454 911 455
rect 901 452 911 454
rect 582 450 588 451
rect 910 451 911 452
rect 915 451 916 455
rect 910 450 916 451
rect 230 446 236 447
rect 766 447 772 448
rect 766 443 767 447
rect 771 446 772 447
rect 858 447 864 448
rect 858 446 859 447
rect 771 444 859 446
rect 771 443 772 444
rect 766 442 772 443
rect 858 443 859 444
rect 863 443 864 447
rect 858 442 864 443
rect 870 447 876 448
rect 870 443 871 447
rect 875 446 876 447
rect 918 447 924 448
rect 918 446 919 447
rect 875 444 919 446
rect 875 443 876 444
rect 870 442 876 443
rect 918 443 919 444
rect 923 443 924 447
rect 918 442 924 443
rect 714 439 720 440
rect 146 435 152 436
rect 146 431 147 435
rect 151 434 152 435
rect 486 435 492 436
rect 486 434 487 435
rect 151 432 487 434
rect 151 431 152 432
rect 146 430 152 431
rect 486 431 487 432
rect 491 431 492 435
rect 714 435 715 439
rect 719 438 720 439
rect 782 439 788 440
rect 719 436 773 438
rect 719 435 720 436
rect 714 434 720 435
rect 782 435 783 439
rect 787 438 788 439
rect 826 439 832 440
rect 826 438 827 439
rect 787 436 827 438
rect 787 435 788 436
rect 782 434 788 435
rect 826 435 827 436
rect 831 438 832 439
rect 874 439 880 440
rect 874 438 875 439
rect 831 436 875 438
rect 831 435 832 436
rect 826 434 832 435
rect 874 435 875 436
rect 879 435 880 439
rect 874 434 880 435
rect 486 430 492 431
rect 698 431 704 432
rect 192 428 402 430
rect 190 427 196 428
rect 190 423 191 427
rect 195 423 196 427
rect 280 425 282 428
rect 400 426 402 428
rect 554 427 560 428
rect 554 426 555 427
rect 400 425 555 426
rect 401 424 555 425
rect 190 422 196 423
rect 554 423 555 424
rect 559 423 560 427
rect 606 427 612 428
rect 606 426 607 427
rect 569 424 607 426
rect 554 422 560 423
rect 606 423 607 424
rect 611 423 612 427
rect 698 427 699 431
rect 703 430 704 431
rect 790 431 796 432
rect 790 430 791 431
rect 703 428 791 430
rect 703 427 704 428
rect 698 426 704 427
rect 712 425 714 428
rect 790 427 791 428
rect 795 427 796 431
rect 822 431 828 432
rect 822 430 823 431
rect 801 428 823 430
rect 790 426 796 427
rect 822 427 823 428
rect 827 427 828 431
rect 822 426 828 427
rect 862 431 868 432
rect 862 427 863 431
rect 867 427 868 431
rect 862 426 868 427
rect 606 422 612 423
rect 790 423 796 424
rect 790 419 791 423
rect 795 419 796 423
rect 222 418 228 419
rect 134 416 140 417
rect 134 412 135 416
rect 139 412 140 416
rect 134 411 140 412
rect 158 416 164 417
rect 158 412 159 416
rect 163 412 164 416
rect 158 411 164 412
rect 182 416 188 417
rect 182 412 183 416
rect 187 412 188 416
rect 222 414 223 418
rect 227 414 228 418
rect 222 413 228 414
rect 342 418 348 419
rect 342 414 343 418
rect 347 414 348 418
rect 510 418 516 419
rect 342 413 348 414
rect 446 416 452 417
rect 182 411 188 412
rect 446 412 447 416
rect 451 412 452 416
rect 446 411 452 412
rect 470 416 476 417
rect 470 412 471 416
rect 475 412 476 416
rect 510 414 511 418
rect 515 414 516 418
rect 654 418 660 419
rect 790 418 796 419
rect 510 413 516 414
rect 614 416 620 417
rect 470 411 476 412
rect 614 412 615 416
rect 619 412 620 416
rect 654 414 655 418
rect 659 414 660 418
rect 654 413 660 414
rect 926 416 932 417
rect 614 411 620 412
rect 926 412 927 416
rect 931 412 932 416
rect 926 411 932 412
rect 110 409 116 410
rect 110 405 111 409
rect 115 405 116 409
rect 958 409 964 410
rect 110 404 116 405
rect 798 405 804 406
rect 234 403 240 404
rect 234 402 235 403
rect 168 400 235 402
rect 151 395 157 396
rect 168 395 170 400
rect 234 399 235 400
rect 239 399 240 403
rect 798 401 799 405
rect 803 401 804 405
rect 958 405 959 409
rect 963 405 964 409
rect 958 404 964 405
rect 798 400 804 401
rect 918 403 924 404
rect 234 398 240 399
rect 918 399 919 403
rect 923 402 924 403
rect 1011 403 1017 404
rect 1011 402 1012 403
rect 923 400 1012 402
rect 923 399 924 400
rect 918 398 924 399
rect 1011 399 1012 400
rect 1016 399 1017 403
rect 1011 398 1017 399
rect 174 395 180 396
rect 151 394 152 395
rect 145 392 152 394
rect 110 391 116 392
rect 110 387 111 391
rect 115 387 116 391
rect 151 391 152 392
rect 156 391 157 395
rect 151 390 157 391
rect 174 391 175 395
rect 179 391 180 395
rect 174 390 180 391
rect 190 395 196 396
rect 190 391 191 395
rect 195 391 196 395
rect 478 395 484 396
rect 190 390 196 391
rect 222 392 228 393
rect 110 386 116 387
rect 158 384 164 385
rect 146 383 152 384
rect 134 382 140 383
rect 134 378 135 382
rect 139 378 140 382
rect 146 379 147 383
rect 151 379 152 383
rect 158 380 159 384
rect 163 380 164 384
rect 176 382 178 390
rect 222 388 223 392
rect 227 388 228 392
rect 206 387 212 388
rect 222 387 228 388
rect 342 392 348 393
rect 342 388 343 392
rect 347 388 348 392
rect 436 392 457 394
rect 342 387 348 388
rect 426 387 432 388
rect 206 386 207 387
rect 196 384 207 386
rect 173 380 178 382
rect 182 382 188 383
rect 158 379 164 380
rect 146 378 152 379
rect 182 378 183 382
rect 187 378 188 382
rect 196 381 198 384
rect 206 383 207 384
rect 211 383 212 387
rect 206 382 212 383
rect 426 383 427 387
rect 431 386 432 387
rect 436 386 438 392
rect 478 391 479 395
rect 483 391 484 395
rect 606 395 612 396
rect 478 390 484 391
rect 510 392 516 393
rect 510 388 511 392
rect 515 388 516 392
rect 606 391 607 395
rect 611 394 612 395
rect 934 395 940 396
rect 611 392 625 394
rect 654 392 660 393
rect 611 391 612 392
rect 606 390 612 391
rect 654 388 655 392
rect 659 388 660 392
rect 510 387 516 388
rect 626 387 632 388
rect 654 387 660 388
rect 798 392 804 393
rect 798 388 799 392
rect 803 388 804 392
rect 934 391 935 395
rect 939 391 940 395
rect 934 390 940 391
rect 958 391 964 392
rect 798 387 804 388
rect 958 387 959 391
rect 963 387 964 391
rect 431 384 438 386
rect 446 384 452 385
rect 470 384 476 385
rect 431 383 432 384
rect 426 382 432 383
rect 446 380 447 384
rect 451 380 452 384
rect 446 379 452 380
rect 458 383 464 384
rect 458 379 459 383
rect 463 379 464 383
rect 470 380 471 384
rect 475 380 476 384
rect 492 384 505 386
rect 614 384 620 385
rect 492 382 494 384
rect 485 380 494 382
rect 614 380 615 384
rect 619 380 620 384
rect 626 383 627 387
rect 631 383 632 387
rect 958 386 964 387
rect 626 382 632 383
rect 470 379 476 380
rect 614 379 620 380
rect 458 378 464 379
rect 134 377 140 378
rect 182 377 188 378
rect 720 374 722 385
rect 926 384 932 385
rect 738 375 744 376
rect 738 374 739 375
rect 720 372 739 374
rect 210 371 216 372
rect 210 367 211 371
rect 215 367 216 371
rect 210 366 216 367
rect 234 371 240 372
rect 234 367 235 371
rect 239 370 240 371
rect 242 371 248 372
rect 242 370 243 371
rect 239 368 243 370
rect 239 367 240 368
rect 234 366 240 367
rect 242 367 243 368
rect 247 370 248 371
rect 278 371 284 372
rect 278 370 279 371
rect 247 368 279 370
rect 247 367 248 368
rect 242 366 248 367
rect 278 367 279 368
rect 283 367 284 371
rect 454 371 460 372
rect 454 370 455 371
rect 405 368 455 370
rect 278 366 284 367
rect 330 367 336 368
rect 194 359 200 360
rect 194 355 195 359
rect 199 358 200 359
rect 224 358 226 365
rect 330 363 331 367
rect 335 363 336 367
rect 454 367 455 368
rect 459 370 460 371
rect 478 371 484 372
rect 478 370 479 371
rect 459 368 479 370
rect 459 367 460 368
rect 454 366 460 367
rect 478 367 479 368
rect 483 367 484 371
rect 478 366 484 367
rect 486 371 492 372
rect 486 367 487 371
rect 491 370 492 371
rect 518 371 524 372
rect 518 370 519 371
rect 491 368 497 370
rect 513 368 519 370
rect 491 367 492 368
rect 486 366 492 367
rect 518 367 519 368
rect 523 367 524 371
rect 594 371 600 372
rect 594 370 595 371
rect 573 368 595 370
rect 518 366 524 367
rect 594 367 595 368
rect 599 367 600 371
rect 686 371 692 372
rect 686 370 687 371
rect 657 368 687 370
rect 594 366 600 367
rect 686 367 687 368
rect 691 367 692 371
rect 738 371 739 372
rect 743 371 744 375
rect 884 374 886 381
rect 926 380 927 384
rect 931 380 932 384
rect 926 379 932 380
rect 936 374 938 381
rect 884 372 938 374
rect 738 370 744 371
rect 686 366 692 367
rect 714 367 720 368
rect 330 362 336 363
rect 344 362 346 365
rect 518 363 524 364
rect 518 362 519 363
rect 344 360 519 362
rect 322 359 328 360
rect 322 358 323 359
rect 199 356 323 358
rect 199 355 200 356
rect 194 354 200 355
rect 322 355 323 356
rect 327 358 328 359
rect 344 358 346 360
rect 518 359 519 360
rect 523 359 524 363
rect 518 358 524 359
rect 644 360 646 365
rect 714 363 715 367
rect 719 363 720 367
rect 714 362 720 363
rect 774 363 780 364
rect 644 359 652 360
rect 327 356 346 358
rect 644 356 647 359
rect 327 355 328 356
rect 322 354 328 355
rect 646 355 647 356
rect 651 355 652 359
rect 774 359 775 363
rect 779 359 780 363
rect 774 358 780 359
rect 834 363 840 364
rect 834 359 835 363
rect 839 362 840 363
rect 839 360 845 362
rect 839 359 840 360
rect 834 358 840 359
rect 646 354 652 355
rect 666 355 672 356
rect 206 351 212 352
rect 206 347 207 351
rect 211 350 212 351
rect 666 351 667 355
rect 671 354 672 355
rect 792 354 794 357
rect 910 355 916 356
rect 910 354 911 355
rect 671 352 911 354
rect 671 351 672 352
rect 666 350 672 351
rect 910 351 911 352
rect 915 351 916 355
rect 910 350 916 351
rect 211 348 334 350
rect 211 347 212 348
rect 206 346 212 347
rect 214 335 220 336
rect 214 331 215 335
rect 219 334 220 335
rect 286 335 292 336
rect 286 334 287 335
rect 219 332 287 334
rect 219 331 220 332
rect 214 330 220 331
rect 286 331 287 332
rect 291 331 292 335
rect 286 330 292 331
rect 298 335 304 336
rect 298 331 299 335
rect 303 331 304 335
rect 322 335 328 336
rect 322 334 323 335
rect 313 332 323 334
rect 298 330 304 331
rect 322 331 323 332
rect 327 331 328 335
rect 332 333 334 348
rect 518 347 524 348
rect 518 343 519 347
rect 523 346 524 347
rect 582 347 588 348
rect 582 346 583 347
rect 523 344 583 346
rect 523 343 524 344
rect 518 342 524 343
rect 582 343 583 344
rect 587 346 588 347
rect 686 347 692 348
rect 686 346 687 347
rect 587 344 687 346
rect 587 343 588 344
rect 582 342 588 343
rect 686 343 687 344
rect 691 343 692 347
rect 862 347 868 348
rect 862 346 863 347
rect 776 344 793 346
rect 800 344 863 346
rect 686 342 692 343
rect 774 343 780 344
rect 658 339 664 340
rect 658 335 659 339
rect 663 338 664 339
rect 698 339 704 340
rect 698 338 699 339
rect 663 336 699 338
rect 663 335 664 336
rect 658 334 664 335
rect 698 335 699 336
rect 703 335 704 339
rect 774 339 775 343
rect 779 339 780 343
rect 774 338 780 339
rect 782 339 788 340
rect 698 334 704 335
rect 782 335 783 339
rect 787 338 788 339
rect 800 338 802 344
rect 862 343 863 344
rect 867 343 868 347
rect 934 347 940 348
rect 934 346 935 347
rect 896 344 935 346
rect 862 342 868 343
rect 874 343 880 344
rect 830 339 836 340
rect 830 338 831 339
rect 787 336 802 338
rect 809 336 831 338
rect 787 335 788 336
rect 782 334 788 335
rect 830 335 831 336
rect 835 335 836 339
rect 874 339 875 343
rect 879 339 880 343
rect 896 342 898 344
rect 934 343 935 344
rect 939 343 940 347
rect 934 342 940 343
rect 893 340 898 342
rect 874 338 880 339
rect 902 339 908 340
rect 830 334 836 335
rect 902 335 903 339
rect 907 335 908 339
rect 902 334 908 335
rect 393 332 411 334
rect 322 330 328 331
rect 409 328 411 332
rect 650 331 656 332
rect 150 327 156 328
rect 150 323 151 327
rect 155 326 156 327
rect 194 327 200 328
rect 194 326 195 327
rect 155 324 169 326
rect 185 324 195 326
rect 155 323 156 324
rect 150 322 156 323
rect 194 323 195 324
rect 199 323 200 327
rect 194 322 200 323
rect 206 327 212 328
rect 206 323 207 327
rect 211 323 212 327
rect 270 327 276 328
rect 270 326 271 327
rect 265 324 271 326
rect 206 322 212 323
rect 270 323 271 324
rect 275 323 276 327
rect 270 322 276 323
rect 407 327 413 328
rect 407 323 408 327
rect 412 326 413 327
rect 490 327 496 328
rect 412 324 481 326
rect 412 323 413 324
rect 407 322 413 323
rect 490 323 491 327
rect 495 323 496 327
rect 490 322 496 323
rect 546 327 552 328
rect 546 323 547 327
rect 551 323 552 327
rect 650 327 651 331
rect 655 330 656 331
rect 742 331 748 332
rect 742 330 743 331
rect 655 328 743 330
rect 655 327 656 328
rect 650 326 656 327
rect 742 327 743 328
rect 747 327 748 331
rect 742 326 748 327
rect 681 324 690 326
rect 546 322 552 323
rect 666 323 672 324
rect 666 319 667 323
rect 671 319 672 323
rect 666 318 672 319
rect 686 323 692 324
rect 686 319 687 323
rect 691 319 692 323
rect 686 318 692 319
rect 698 323 704 324
rect 698 319 699 323
rect 703 319 704 323
rect 862 323 868 324
rect 862 322 863 323
rect 733 320 863 322
rect 698 318 704 319
rect 862 319 863 320
rect 867 319 868 323
rect 862 318 868 319
rect 742 315 748 316
rect 286 311 292 312
rect 286 307 287 311
rect 291 310 292 311
rect 334 311 340 312
rect 334 310 335 311
rect 291 308 335 310
rect 291 307 292 308
rect 286 306 292 307
rect 334 307 335 308
rect 339 307 340 311
rect 742 311 743 315
rect 747 314 748 315
rect 902 315 908 316
rect 902 314 903 315
rect 747 312 858 314
rect 747 311 748 312
rect 742 310 748 311
rect 856 310 858 312
rect 872 312 903 314
rect 872 310 874 312
rect 902 311 903 312
rect 907 311 908 315
rect 902 310 908 311
rect 918 311 924 312
rect 856 308 874 310
rect 650 307 656 308
rect 334 306 340 307
rect 414 306 420 307
rect 134 304 140 305
rect 134 300 135 304
rect 139 300 140 304
rect 158 303 164 304
rect 158 302 159 303
rect 149 300 159 302
rect 134 299 140 300
rect 158 299 159 300
rect 163 299 164 303
rect 414 302 415 306
rect 419 302 420 306
rect 638 306 644 307
rect 438 304 444 305
rect 414 301 420 302
rect 426 303 432 304
rect 158 298 164 299
rect 426 299 427 303
rect 431 299 432 303
rect 438 300 439 304
rect 443 300 444 304
rect 638 302 639 306
rect 643 302 644 306
rect 650 303 651 307
rect 655 303 656 307
rect 766 307 772 308
rect 766 306 767 307
rect 745 304 767 306
rect 650 302 656 303
rect 766 303 767 304
rect 771 303 772 307
rect 766 302 772 303
rect 878 307 884 308
rect 878 303 879 307
rect 883 303 884 307
rect 918 307 919 311
rect 923 310 924 311
rect 923 308 938 310
rect 923 307 924 308
rect 918 306 924 307
rect 878 302 884 303
rect 926 304 932 305
rect 453 300 489 302
rect 638 301 644 302
rect 926 300 927 304
rect 931 300 932 304
rect 936 301 938 308
rect 438 299 444 300
rect 926 299 932 300
rect 426 298 432 299
rect 110 297 116 298
rect 958 297 964 298
rect 110 293 111 297
rect 115 293 116 297
rect 110 292 116 293
rect 182 296 188 297
rect 182 292 183 296
rect 187 292 188 296
rect 182 291 188 292
rect 310 296 316 297
rect 310 292 311 296
rect 315 292 316 296
rect 502 296 508 297
rect 678 296 684 297
rect 502 292 503 296
rect 507 292 508 296
rect 658 295 664 296
rect 658 294 659 295
rect 649 292 659 294
rect 310 291 316 292
rect 407 291 413 292
rect 144 286 146 289
rect 206 287 212 288
rect 206 286 207 287
rect 144 284 207 286
rect 206 283 207 284
rect 211 283 212 287
rect 407 287 408 291
rect 412 290 413 291
rect 422 291 428 292
rect 422 290 423 291
rect 412 288 423 290
rect 412 287 413 288
rect 407 286 413 287
rect 422 287 423 288
rect 427 287 428 291
rect 494 291 500 292
rect 502 291 508 292
rect 658 291 659 292
rect 663 291 664 295
rect 678 292 679 296
rect 683 292 684 296
rect 678 291 684 292
rect 806 295 812 296
rect 806 291 807 295
rect 811 291 812 295
rect 958 293 959 297
rect 963 293 964 297
rect 958 292 964 293
rect 494 290 495 291
rect 449 289 495 290
rect 422 286 428 287
rect 448 288 495 289
rect 448 284 450 288
rect 494 287 495 288
rect 499 287 500 291
rect 658 290 664 291
rect 806 290 812 291
rect 862 291 868 292
rect 494 286 500 287
rect 862 287 863 291
rect 867 290 868 291
rect 946 291 952 292
rect 946 290 947 291
rect 867 288 947 290
rect 867 287 868 288
rect 862 286 868 287
rect 946 287 947 288
rect 951 287 952 291
rect 946 286 952 287
rect 206 282 212 283
rect 446 283 452 284
rect 110 279 116 280
rect 110 275 111 279
rect 115 275 116 279
rect 110 274 116 275
rect 310 279 316 280
rect 310 275 311 279
rect 315 275 316 279
rect 446 279 447 283
rect 451 279 452 283
rect 446 278 452 279
rect 502 283 508 284
rect 502 279 503 283
rect 507 279 508 283
rect 502 278 508 279
rect 678 282 684 283
rect 678 278 679 282
rect 683 278 684 282
rect 958 279 964 280
rect 678 277 684 278
rect 802 277 808 278
rect 310 274 316 275
rect 802 273 803 277
rect 807 273 808 277
rect 958 275 959 279
rect 963 275 964 279
rect 958 274 964 275
rect 134 272 140 273
rect 134 268 135 272
rect 139 268 140 272
rect 134 267 140 268
rect 198 272 204 273
rect 198 268 199 272
rect 203 268 204 272
rect 414 272 420 273
rect 414 268 415 272
rect 419 268 420 272
rect 198 267 204 268
rect 346 267 352 268
rect 414 267 420 268
rect 438 272 444 273
rect 638 272 644 273
rect 802 272 808 273
rect 926 272 932 273
rect 438 268 439 272
rect 443 268 444 272
rect 438 267 444 268
rect 447 271 453 272
rect 447 267 448 271
rect 452 270 453 271
rect 486 271 492 272
rect 486 270 487 271
rect 452 268 487 270
rect 452 267 453 268
rect 346 266 347 267
rect 184 260 186 265
rect 317 264 347 266
rect 346 263 347 264
rect 351 263 352 267
rect 447 266 453 267
rect 486 267 487 268
rect 491 267 492 271
rect 638 268 639 272
rect 643 268 644 272
rect 638 267 644 268
rect 926 268 927 272
rect 931 268 932 272
rect 926 267 932 268
rect 486 266 492 267
rect 346 262 352 263
rect 554 263 560 264
rect 158 259 164 260
rect 158 255 159 259
rect 163 255 164 259
rect 158 254 164 255
rect 174 259 180 260
rect 174 255 175 259
rect 179 255 180 259
rect 174 254 180 255
rect 182 259 188 260
rect 182 255 183 259
rect 187 255 188 259
rect 294 259 300 260
rect 182 254 188 255
rect 242 255 248 256
rect 242 251 243 255
rect 247 251 248 255
rect 294 255 295 259
rect 299 255 300 259
rect 294 254 300 255
rect 318 259 324 260
rect 318 255 319 259
rect 323 258 324 259
rect 554 259 555 263
rect 559 262 560 263
rect 646 263 652 264
rect 646 262 647 263
rect 559 260 647 262
rect 559 259 560 260
rect 554 258 560 259
rect 646 259 647 260
rect 651 259 652 263
rect 646 258 652 259
rect 774 259 780 260
rect 323 256 377 258
rect 323 255 324 256
rect 318 254 324 255
rect 462 255 468 256
rect 462 254 463 255
rect 242 250 248 251
rect 158 247 164 248
rect 158 243 159 247
rect 163 246 164 247
rect 296 246 298 254
rect 449 252 463 254
rect 302 251 308 252
rect 302 247 303 251
rect 307 250 308 251
rect 449 250 451 252
rect 462 251 463 252
rect 467 251 468 255
rect 566 255 572 256
rect 462 250 468 251
rect 307 248 451 250
rect 307 247 308 248
rect 302 246 308 247
rect 454 247 461 248
rect 163 244 298 246
rect 163 243 164 244
rect 158 242 164 243
rect 454 243 455 247
rect 460 246 461 247
rect 486 247 492 248
rect 460 244 477 246
rect 460 243 461 244
rect 454 242 461 243
rect 486 243 487 247
rect 491 243 492 247
rect 504 246 506 253
rect 566 251 567 255
rect 571 251 572 255
rect 774 255 775 259
rect 779 258 780 259
rect 934 259 940 260
rect 934 258 935 259
rect 779 256 935 258
rect 779 255 780 256
rect 774 254 780 255
rect 934 255 935 256
rect 939 255 940 259
rect 934 254 940 255
rect 566 250 572 251
rect 742 247 748 248
rect 742 246 743 247
rect 504 244 743 246
rect 486 242 492 243
rect 742 243 743 244
rect 747 243 748 247
rect 742 242 748 243
rect 284 240 442 242
rect 158 239 164 240
rect 158 235 159 239
rect 163 238 164 239
rect 242 239 248 240
rect 242 238 243 239
rect 163 236 243 238
rect 163 235 164 236
rect 158 234 164 235
rect 242 235 243 236
rect 247 235 248 239
rect 242 234 248 235
rect 206 231 212 232
rect 206 227 207 231
rect 211 230 212 231
rect 238 231 244 232
rect 284 231 286 240
rect 390 235 396 236
rect 390 234 391 235
rect 333 232 391 234
rect 390 231 391 232
rect 395 231 396 235
rect 440 232 442 240
rect 466 235 472 236
rect 238 230 239 231
rect 211 228 239 230
rect 211 227 212 228
rect 206 226 212 227
rect 238 227 239 228
rect 243 227 244 231
rect 390 230 396 231
rect 438 231 444 232
rect 238 226 244 227
rect 438 227 439 231
rect 443 227 444 231
rect 466 231 467 235
rect 471 234 472 235
rect 566 235 572 236
rect 566 234 567 235
rect 471 232 567 234
rect 471 231 472 232
rect 466 230 472 231
rect 566 231 567 232
rect 571 231 572 235
rect 566 230 572 231
rect 438 226 444 227
rect 142 224 148 225
rect 142 220 143 224
rect 147 220 148 224
rect 142 219 148 220
rect 166 224 172 225
rect 166 220 167 224
rect 171 220 172 224
rect 166 219 172 220
rect 190 224 196 225
rect 382 224 388 225
rect 190 220 191 224
rect 195 220 196 224
rect 190 219 196 220
rect 278 223 284 224
rect 278 219 279 223
rect 283 219 284 223
rect 382 220 383 224
rect 387 220 388 224
rect 382 219 388 220
rect 406 224 412 225
rect 406 220 407 224
rect 411 220 412 224
rect 406 219 412 220
rect 430 224 436 225
rect 430 220 431 224
rect 435 220 436 224
rect 734 224 740 225
rect 734 220 735 224
rect 739 220 740 224
rect 430 219 436 220
rect 474 219 480 220
rect 734 219 740 220
rect 774 224 780 225
rect 774 220 775 224
rect 779 220 780 224
rect 774 219 780 220
rect 814 224 820 225
rect 814 220 815 224
rect 819 220 820 224
rect 814 219 820 220
rect 854 224 860 225
rect 854 220 855 224
rect 859 220 860 224
rect 854 219 860 220
rect 902 224 908 225
rect 902 220 903 224
rect 907 220 908 224
rect 902 219 908 220
rect 926 224 932 225
rect 926 220 927 224
rect 931 220 932 224
rect 926 219 932 220
rect 278 218 284 219
rect 110 217 116 218
rect 110 213 111 217
rect 115 213 116 217
rect 474 215 475 219
rect 479 215 480 219
rect 958 217 964 218
rect 474 214 480 215
rect 622 214 628 215
rect 110 212 116 213
rect 390 211 396 212
rect 390 207 391 211
rect 395 210 396 211
rect 446 211 453 212
rect 446 210 447 211
rect 395 208 447 210
rect 395 207 396 208
rect 390 206 396 207
rect 446 207 447 208
rect 452 207 453 211
rect 622 210 623 214
rect 627 210 628 214
rect 958 213 959 217
rect 963 213 964 217
rect 958 212 964 213
rect 622 209 628 210
rect 446 206 453 207
rect 534 207 540 208
rect 135 203 141 204
rect 110 199 116 200
rect 110 195 111 199
rect 115 195 116 199
rect 135 199 136 203
rect 140 202 141 203
rect 150 203 156 204
rect 150 202 151 203
rect 140 200 151 202
rect 140 199 141 200
rect 135 198 141 199
rect 150 199 151 200
rect 155 199 156 203
rect 190 203 196 204
rect 392 203 394 206
rect 454 203 460 204
rect 190 202 191 203
rect 177 200 191 202
rect 150 198 156 199
rect 190 199 191 200
rect 195 199 196 203
rect 454 202 455 203
rect 201 200 214 202
rect 190 198 196 199
rect 110 194 116 195
rect 154 195 160 196
rect 142 192 148 193
rect 142 188 143 192
rect 147 188 148 192
rect 154 191 155 195
rect 159 191 160 195
rect 178 195 184 196
rect 154 190 160 191
rect 166 192 172 193
rect 142 187 148 188
rect 166 188 167 192
rect 171 188 172 192
rect 178 191 179 195
rect 183 191 184 195
rect 178 190 184 191
rect 190 192 196 193
rect 166 187 172 188
rect 190 188 191 192
rect 195 188 196 192
rect 190 187 196 188
rect 202 191 208 192
rect 202 187 203 191
rect 207 187 208 191
rect 212 188 214 200
rect 400 200 417 202
rect 441 200 455 202
rect 302 195 308 196
rect 302 191 303 195
rect 307 191 308 195
rect 302 190 308 191
rect 382 192 388 193
rect 400 192 402 200
rect 454 199 455 200
rect 459 202 460 203
rect 466 203 472 204
rect 466 202 467 203
rect 459 200 467 202
rect 459 199 460 200
rect 454 198 460 199
rect 466 199 467 200
rect 471 199 472 203
rect 534 203 535 207
rect 539 206 540 207
rect 591 207 597 208
rect 591 206 592 207
rect 539 204 592 206
rect 539 203 540 204
rect 534 202 540 203
rect 591 203 592 204
rect 596 203 597 207
rect 591 202 597 203
rect 742 203 748 204
rect 466 198 472 199
rect 474 200 480 201
rect 474 196 475 200
rect 479 196 480 200
rect 474 195 480 196
rect 622 200 628 201
rect 622 196 623 200
rect 627 196 628 200
rect 742 199 743 203
rect 747 199 748 203
rect 742 198 748 199
rect 782 203 788 204
rect 782 199 783 203
rect 787 199 788 203
rect 782 198 788 199
rect 822 203 828 204
rect 822 199 823 203
rect 827 199 828 203
rect 886 203 892 204
rect 886 202 887 203
rect 865 200 887 202
rect 822 198 828 199
rect 886 199 887 200
rect 891 199 892 203
rect 886 198 892 199
rect 910 203 916 204
rect 910 199 911 203
rect 915 199 916 203
rect 910 198 916 199
rect 934 203 940 204
rect 934 199 935 203
rect 939 199 940 203
rect 934 198 940 199
rect 958 199 964 200
rect 622 195 628 196
rect 958 195 959 199
rect 963 195 964 199
rect 958 194 964 195
rect 382 188 383 192
rect 387 188 388 192
rect 202 186 208 187
rect 210 187 216 188
rect 210 183 211 187
rect 215 183 216 187
rect 210 182 216 183
rect 218 187 224 188
rect 382 187 388 188
rect 394 191 402 192
rect 394 187 395 191
rect 399 188 402 191
rect 406 192 412 193
rect 406 188 407 192
rect 411 188 412 192
rect 430 192 436 193
rect 734 192 740 193
rect 774 192 780 193
rect 421 188 426 190
rect 399 187 400 188
rect 406 187 412 188
rect 218 183 219 187
rect 223 183 224 187
rect 394 186 400 187
rect 218 182 224 183
rect 424 182 426 188
rect 430 188 431 192
rect 435 188 436 192
rect 455 191 461 192
rect 455 190 456 191
rect 445 188 456 190
rect 430 187 436 188
rect 455 187 456 188
rect 460 187 461 191
rect 634 191 640 192
rect 455 186 461 187
rect 468 182 470 189
rect 634 187 635 191
rect 639 187 640 191
rect 734 188 735 192
rect 739 188 740 192
rect 734 187 740 188
rect 746 191 752 192
rect 746 187 747 191
rect 751 187 752 191
rect 774 188 775 192
rect 779 188 780 192
rect 814 192 820 193
rect 774 187 780 188
rect 634 186 640 187
rect 746 186 752 187
rect 424 180 470 182
rect 574 183 580 184
rect 135 179 141 180
rect 135 175 136 179
rect 140 178 141 179
rect 574 179 575 183
rect 579 182 580 183
rect 598 183 604 184
rect 598 182 599 183
rect 579 180 599 182
rect 579 179 580 180
rect 574 178 580 179
rect 598 179 599 180
rect 603 179 604 183
rect 598 178 604 179
rect 714 183 720 184
rect 714 179 715 183
rect 719 182 720 183
rect 758 183 764 184
rect 758 182 759 183
rect 719 180 759 182
rect 719 179 720 180
rect 714 178 720 179
rect 758 179 759 180
rect 763 182 764 183
rect 784 182 786 189
rect 814 188 815 192
rect 819 188 820 192
rect 854 192 860 193
rect 902 192 908 193
rect 814 187 820 188
rect 763 180 786 182
rect 824 182 826 189
rect 854 188 855 192
rect 859 188 860 192
rect 878 191 884 192
rect 878 190 879 191
rect 869 188 879 190
rect 854 187 860 188
rect 878 187 879 188
rect 883 187 884 191
rect 902 188 903 192
rect 907 188 908 192
rect 946 191 952 192
rect 926 190 932 191
rect 946 190 947 191
rect 902 187 908 188
rect 878 186 884 187
rect 830 183 836 184
rect 830 182 831 183
rect 824 180 831 182
rect 763 179 764 180
rect 758 178 764 179
rect 140 176 234 178
rect 140 175 141 176
rect 135 174 141 175
rect 232 170 234 176
rect 262 177 268 178
rect 262 173 263 177
rect 267 173 268 177
rect 368 176 578 178
rect 368 174 370 176
rect 746 175 752 176
rect 262 172 268 173
rect 337 172 370 174
rect 460 172 610 174
rect 318 171 324 172
rect 318 170 319 171
rect 232 168 319 170
rect 318 167 319 168
rect 323 167 324 171
rect 318 166 324 167
rect 334 171 342 172
rect 334 167 335 171
rect 339 168 342 171
rect 446 171 452 172
rect 339 167 340 168
rect 334 166 340 167
rect 446 167 447 171
rect 451 170 452 171
rect 460 170 462 172
rect 451 168 462 170
rect 608 169 610 172
rect 631 171 637 172
rect 631 170 632 171
rect 625 168 632 170
rect 451 167 452 168
rect 446 166 452 167
rect 631 167 632 168
rect 636 167 637 171
rect 631 166 637 167
rect 642 171 648 172
rect 642 167 643 171
rect 647 167 648 171
rect 746 171 747 175
rect 751 174 752 175
rect 824 174 826 180
rect 830 179 831 180
rect 835 179 836 183
rect 830 178 836 179
rect 886 183 892 184
rect 886 179 887 183
rect 891 182 892 183
rect 912 182 914 189
rect 926 186 927 190
rect 931 186 932 190
rect 941 188 947 190
rect 946 187 947 188
rect 951 187 952 191
rect 946 186 952 187
rect 926 185 932 186
rect 891 180 914 182
rect 891 179 892 180
rect 886 178 892 179
rect 751 172 826 174
rect 751 171 752 172
rect 746 170 752 171
rect 642 166 648 167
rect 202 163 208 164
rect 202 159 203 163
rect 207 162 208 163
rect 270 163 276 164
rect 207 160 261 162
rect 207 159 208 160
rect 202 158 208 159
rect 270 159 271 163
rect 275 162 276 163
rect 326 163 332 164
rect 326 162 327 163
rect 275 160 281 162
rect 309 160 327 162
rect 275 159 276 160
rect 270 158 276 159
rect 326 159 327 160
rect 331 159 332 163
rect 326 158 332 159
rect 591 163 597 164
rect 591 159 592 163
rect 596 162 597 163
rect 676 162 678 167
rect 596 160 678 162
rect 596 159 597 160
rect 591 158 597 159
rect 454 155 460 156
rect 454 151 455 155
rect 459 151 460 155
rect 486 155 492 156
rect 454 150 460 151
rect 481 148 483 154
rect 486 151 487 155
rect 491 154 492 155
rect 574 155 580 156
rect 491 152 549 154
rect 491 151 492 152
rect 486 150 492 151
rect 238 147 244 148
rect 238 143 239 147
rect 243 143 244 147
rect 270 147 276 148
rect 270 143 271 147
rect 275 146 276 147
rect 394 147 400 148
rect 394 146 395 147
rect 275 144 395 146
rect 275 143 276 144
rect 238 142 244 143
rect 210 139 216 140
rect 210 135 211 139
rect 215 138 216 139
rect 252 138 254 143
rect 270 142 276 143
rect 394 143 395 144
rect 399 143 400 147
rect 479 147 485 148
rect 394 142 400 143
rect 422 143 428 144
rect 319 140 390 142
rect 319 138 321 140
rect 215 136 321 138
rect 215 135 216 136
rect 210 134 216 135
rect 346 135 352 136
rect 346 131 347 135
rect 351 134 352 135
rect 388 134 390 140
rect 422 139 423 143
rect 427 142 428 143
rect 468 142 470 145
rect 479 143 480 147
rect 484 143 485 147
rect 479 142 485 143
rect 494 147 500 148
rect 494 143 495 147
rect 499 146 500 147
rect 560 146 562 153
rect 574 151 575 155
rect 579 151 580 155
rect 574 150 580 151
rect 631 155 637 156
rect 631 151 632 155
rect 636 154 637 155
rect 686 155 692 156
rect 686 154 687 155
rect 636 152 687 154
rect 636 151 637 152
rect 631 150 637 151
rect 686 151 687 152
rect 691 154 692 155
rect 746 155 752 156
rect 746 154 747 155
rect 691 152 747 154
rect 691 151 692 152
rect 686 150 692 151
rect 746 151 747 152
rect 751 151 752 155
rect 746 150 752 151
rect 499 144 562 146
rect 499 143 500 144
rect 494 142 500 143
rect 631 143 637 144
rect 631 142 632 143
rect 427 140 470 142
rect 504 140 632 142
rect 427 139 428 140
rect 422 138 428 139
rect 495 139 501 140
rect 486 135 492 136
rect 486 134 487 135
rect 351 132 378 134
rect 388 132 487 134
rect 351 131 352 132
rect 346 130 352 131
rect 134 128 140 129
rect 134 124 135 128
rect 139 124 140 128
rect 238 128 244 129
rect 149 124 230 126
rect 134 123 140 124
rect 110 121 116 122
rect 110 117 111 121
rect 115 117 116 121
rect 218 119 224 120
rect 218 118 219 119
rect 110 116 116 117
rect 145 116 219 118
rect 218 115 219 116
rect 223 115 224 119
rect 228 118 230 124
rect 238 124 239 128
rect 243 124 244 128
rect 366 128 372 129
rect 253 124 321 126
rect 238 123 244 124
rect 319 118 321 124
rect 366 124 367 128
rect 371 124 372 128
rect 376 125 378 132
rect 486 131 487 132
rect 491 131 492 135
rect 495 135 496 139
rect 500 138 501 139
rect 504 138 506 140
rect 631 139 632 140
rect 636 139 637 143
rect 631 138 637 139
rect 500 136 506 138
rect 500 135 501 136
rect 495 134 501 135
rect 551 135 557 136
rect 486 130 492 131
rect 551 131 552 135
rect 556 134 557 135
rect 556 132 762 134
rect 556 131 557 132
rect 551 130 557 131
rect 494 128 500 129
rect 366 123 372 124
rect 494 124 495 128
rect 499 124 500 128
rect 622 128 628 129
rect 750 128 756 129
rect 494 123 500 124
rect 508 122 510 125
rect 622 124 623 128
rect 627 124 628 128
rect 622 123 628 124
rect 634 127 640 128
rect 634 123 635 127
rect 639 123 640 127
rect 750 124 751 128
rect 755 124 756 128
rect 760 125 762 132
rect 750 123 756 124
rect 634 122 640 123
rect 508 120 606 122
rect 604 118 606 120
rect 958 121 964 122
rect 228 116 249 118
rect 319 116 377 118
rect 604 116 633 118
rect 958 117 959 121
rect 963 117 964 121
rect 958 116 964 117
rect 218 114 224 115
rect 438 115 444 116
rect 438 111 439 115
rect 443 114 444 115
rect 546 115 552 116
rect 546 114 547 115
rect 443 112 547 114
rect 443 111 444 112
rect 438 110 444 111
rect 546 111 547 112
rect 551 111 552 115
rect 546 110 552 111
rect 758 115 764 116
rect 758 111 759 115
rect 763 111 764 115
rect 758 110 764 111
rect 110 103 116 104
rect 110 99 111 103
rect 115 99 116 103
rect 110 98 116 99
rect 958 103 964 104
rect 958 99 959 103
rect 963 99 964 103
rect 958 98 964 99
rect 134 96 140 97
rect 134 92 135 96
rect 139 92 140 96
rect 134 91 140 92
rect 238 96 244 97
rect 238 92 239 96
rect 243 92 244 96
rect 238 91 244 92
rect 366 96 372 97
rect 366 92 367 96
rect 371 92 372 96
rect 366 91 372 92
rect 494 96 500 97
rect 494 92 495 96
rect 499 92 500 96
rect 494 91 500 92
rect 622 96 628 97
rect 622 92 623 96
rect 627 92 628 96
rect 622 91 628 92
rect 750 96 756 97
rect 750 92 751 96
rect 755 92 756 96
rect 750 91 756 92
<< m3c >>
rect 135 996 139 1000
rect 319 996 323 1000
rect 527 996 531 1000
rect 735 996 739 1000
rect 927 996 931 1000
rect 111 989 115 993
rect 835 991 839 995
rect 959 989 963 993
rect 939 983 943 987
rect 111 971 115 975
rect 203 975 207 979
rect 135 964 139 968
rect 319 964 323 968
rect 947 975 951 979
rect 527 964 531 968
rect 287 947 291 951
rect 299 947 303 951
rect 319 947 323 951
rect 427 955 431 959
rect 735 964 739 968
rect 759 963 763 967
rect 927 964 931 968
rect 939 967 943 971
rect 959 971 963 975
rect 443 947 447 951
rect 299 923 303 927
rect 135 916 139 920
rect 147 915 151 919
rect 159 916 163 920
rect 171 915 175 919
rect 183 916 187 920
rect 223 915 227 919
rect 231 916 235 920
rect 251 915 255 919
rect 299 915 303 919
rect 455 916 459 920
rect 467 915 471 919
rect 519 916 523 920
rect 531 915 535 919
rect 583 916 587 920
rect 631 915 635 919
rect 647 916 651 920
rect 667 915 671 919
rect 711 916 715 920
rect 723 915 727 919
rect 111 909 115 913
rect 311 908 315 912
rect 191 903 195 907
rect 371 907 375 911
rect 239 903 243 907
rect 767 916 771 920
rect 815 915 819 919
rect 823 916 827 920
rect 835 915 839 919
rect 887 916 891 920
rect 919 915 923 919
rect 927 916 931 920
rect 947 915 951 919
rect 959 909 963 913
rect 111 891 115 895
rect 251 895 255 899
rect 379 899 383 903
rect 511 899 515 903
rect 539 903 543 907
rect 655 903 659 907
rect 703 903 707 907
rect 843 903 847 907
rect 311 891 315 895
rect 531 891 535 895
rect 835 895 839 899
rect 947 903 951 907
rect 959 891 963 895
rect 135 884 139 888
rect 159 884 163 888
rect 183 884 187 888
rect 231 884 235 888
rect 459 884 463 888
rect 519 884 523 888
rect 583 884 587 888
rect 647 884 651 888
rect 711 884 715 888
rect 767 884 771 888
rect 823 884 827 888
rect 887 884 891 888
rect 927 884 931 888
rect 127 875 131 879
rect 191 875 195 879
rect 275 875 279 879
rect 427 879 431 883
rect 339 871 343 875
rect 347 871 351 875
rect 435 875 439 879
rect 703 875 707 879
rect 147 859 151 863
rect 727 867 731 871
rect 151 851 155 855
rect 223 851 227 855
rect 231 851 235 855
rect 339 855 343 859
rect 539 859 543 863
rect 167 843 171 847
rect 359 843 363 847
rect 379 847 383 851
rect 387 847 391 851
rect 519 847 523 851
rect 527 851 531 855
rect 655 851 659 855
rect 703 851 707 855
rect 727 855 731 859
rect 767 855 771 859
rect 563 843 567 847
rect 899 847 903 851
rect 175 836 179 840
rect 327 835 331 839
rect 575 836 579 840
rect 775 836 779 840
rect 807 836 811 840
rect 847 838 851 842
rect 111 829 115 833
rect 451 831 455 835
rect 275 823 279 827
rect 347 823 351 827
rect 519 827 523 831
rect 587 823 591 827
rect 639 825 643 829
rect 959 829 963 833
rect 111 811 115 815
rect 159 812 163 816
rect 451 812 455 816
rect 595 815 599 819
rect 639 812 643 816
rect 767 815 771 819
rect 847 812 851 816
rect 203 803 207 807
rect 383 799 387 803
rect 471 803 475 807
rect 575 804 579 808
rect 587 807 591 811
rect 959 811 963 815
rect 631 807 635 811
rect 775 804 779 808
rect 275 791 279 795
rect 311 789 315 793
rect 555 795 559 799
rect 739 795 743 799
rect 807 804 811 808
rect 819 803 823 807
rect 827 807 831 811
rect 835 791 839 795
rect 855 791 859 795
rect 127 783 131 787
rect 199 775 203 779
rect 367 783 371 787
rect 375 783 379 787
rect 443 783 447 787
rect 487 783 491 787
rect 299 775 303 779
rect 367 775 371 779
rect 627 779 631 783
rect 431 767 435 771
rect 319 759 323 763
rect 239 751 243 755
rect 367 759 371 763
rect 443 763 447 767
rect 527 767 531 771
rect 539 767 543 771
rect 555 767 559 771
rect 683 767 687 771
rect 511 759 515 763
rect 627 759 631 763
rect 819 759 823 763
rect 527 751 531 755
rect 551 751 555 755
rect 667 751 671 755
rect 711 751 715 755
rect 359 743 363 747
rect 451 743 455 747
rect 479 743 483 747
rect 295 735 299 739
rect 375 735 379 739
rect 507 739 511 743
rect 791 743 795 747
rect 823 743 827 747
rect 835 747 839 751
rect 859 743 860 747
rect 860 743 863 747
rect 867 743 871 747
rect 927 743 931 747
rect 199 727 203 731
rect 231 727 235 731
rect 515 731 519 735
rect 551 731 555 735
rect 563 731 567 735
rect 595 735 599 739
rect 683 735 687 739
rect 711 727 715 731
rect 767 727 771 731
rect 315 719 319 723
rect 135 712 139 716
rect 279 712 283 716
rect 291 711 295 715
rect 303 712 307 716
rect 327 712 331 716
rect 339 711 343 715
rect 351 714 355 718
rect 375 715 379 719
rect 383 712 387 716
rect 407 711 411 715
rect 415 714 419 718
rect 439 712 443 716
rect 451 711 455 715
rect 463 712 467 716
rect 495 714 499 718
rect 507 715 511 719
rect 919 719 923 723
rect 655 712 659 716
rect 799 712 803 716
rect 835 711 839 715
rect 111 705 115 709
rect 175 704 179 708
rect 143 699 147 703
rect 287 699 291 703
rect 111 687 115 691
rect 359 699 363 703
rect 391 699 395 703
rect 423 699 427 703
rect 447 699 451 703
rect 487 703 491 707
rect 543 704 547 708
rect 695 704 699 708
rect 847 704 851 708
rect 959 705 963 709
rect 407 691 411 695
rect 487 695 491 699
rect 663 699 667 703
rect 807 699 811 703
rect 543 690 547 694
rect 847 687 851 691
rect 959 687 963 691
rect 135 680 139 684
rect 175 678 179 682
rect 279 680 283 684
rect 303 680 307 684
rect 327 680 331 684
rect 351 680 355 684
rect 383 680 387 684
rect 415 680 419 684
rect 439 680 443 684
rect 463 680 467 684
rect 495 680 499 684
rect 655 680 659 684
rect 695 678 699 682
rect 799 680 803 684
rect 151 671 155 675
rect 359 671 363 675
rect 563 671 567 675
rect 759 671 763 675
rect 143 663 147 667
rect 319 663 323 667
rect 671 663 675 667
rect 835 667 839 671
rect 939 675 943 679
rect 295 647 299 651
rect 275 639 279 643
rect 467 643 471 647
rect 595 647 599 651
rect 663 655 667 659
rect 807 659 811 663
rect 819 659 823 663
rect 263 627 267 631
rect 335 631 339 635
rect 431 631 435 635
rect 567 635 571 639
rect 619 639 623 643
rect 639 647 643 651
rect 679 639 683 643
rect 831 647 835 651
rect 811 639 815 643
rect 607 631 611 635
rect 303 624 307 628
rect 455 623 459 627
rect 559 624 563 628
rect 583 624 587 628
rect 775 624 779 628
rect 799 627 803 631
rect 839 624 843 628
rect 927 624 931 628
rect 111 617 115 621
rect 159 617 163 621
rect 231 607 235 611
rect 275 607 279 611
rect 359 607 363 611
rect 511 611 515 615
rect 539 611 543 615
rect 647 613 651 617
rect 959 617 963 621
rect 111 599 115 603
rect 159 600 163 604
rect 287 600 291 604
rect 551 603 555 607
rect 567 603 571 607
rect 639 603 643 607
rect 647 600 651 604
rect 783 603 787 607
rect 823 600 827 604
rect 199 587 203 591
rect 279 587 283 591
rect 327 591 331 595
rect 479 595 483 599
rect 559 592 563 596
rect 571 591 575 595
rect 583 592 587 596
rect 595 591 599 595
rect 775 592 779 596
rect 383 579 387 583
rect 799 591 803 595
rect 867 595 871 599
rect 959 599 963 603
rect 927 592 931 596
rect 939 591 943 595
rect 791 583 792 587
rect 792 583 795 587
rect 439 577 443 581
rect 135 559 139 563
rect 147 559 151 563
rect 239 559 243 563
rect 279 567 283 571
rect 295 571 296 575
rect 296 571 299 575
rect 351 571 355 575
rect 383 559 387 563
rect 411 563 415 567
rect 671 571 675 575
rect 795 571 799 575
rect 815 571 819 575
rect 455 563 459 567
rect 831 567 835 571
rect 847 571 851 575
rect 867 571 871 575
rect 879 567 883 571
rect 483 555 487 559
rect 551 559 555 563
rect 811 559 815 563
rect 947 559 951 563
rect 455 547 459 551
rect 571 551 575 555
rect 711 551 715 555
rect 831 551 835 555
rect 871 551 875 555
rect 239 539 243 543
rect 359 531 363 535
rect 371 535 375 539
rect 391 535 395 539
rect 615 535 619 539
rect 847 543 851 547
rect 439 527 443 531
rect 467 527 471 531
rect 483 527 487 531
rect 839 535 843 539
rect 491 523 495 527
rect 143 515 147 519
rect 139 507 143 511
rect 551 515 555 519
rect 583 515 587 519
rect 607 515 611 519
rect 763 519 767 523
rect 783 523 787 527
rect 907 527 911 531
rect 871 519 875 523
rect 371 507 375 511
rect 423 507 427 511
rect 795 507 799 511
rect 311 499 315 503
rect 687 499 691 503
rect 711 499 715 503
rect 811 503 815 507
rect 831 507 835 511
rect 879 511 883 515
rect 175 491 179 495
rect 255 492 259 496
rect 267 491 271 495
rect 279 492 283 496
rect 291 491 295 495
rect 303 492 307 496
rect 327 492 331 496
rect 519 492 523 496
rect 627 491 631 495
rect 703 492 707 496
rect 751 492 755 496
rect 763 491 767 495
rect 871 495 875 499
rect 111 485 115 489
rect 151 484 155 488
rect 279 479 283 483
rect 303 479 307 483
rect 319 483 323 487
rect 351 483 355 487
rect 379 484 383 488
rect 431 483 435 487
rect 459 483 463 487
rect 467 483 471 487
rect 575 484 579 488
rect 679 483 683 487
rect 959 485 963 489
rect 447 475 451 479
rect 491 475 495 479
rect 111 467 115 471
rect 575 470 579 474
rect 783 471 787 475
rect 379 465 383 469
rect 151 458 155 462
rect 255 460 259 464
rect 279 460 283 464
rect 303 460 307 464
rect 327 460 331 464
rect 519 460 523 464
rect 703 460 707 464
rect 751 460 755 464
rect 775 463 779 467
rect 911 475 915 479
rect 959 467 963 471
rect 847 461 851 465
rect 231 447 235 451
rect 439 451 443 455
rect 583 451 587 455
rect 763 455 767 459
rect 835 455 839 459
rect 911 451 915 455
rect 767 443 771 447
rect 859 443 863 447
rect 871 443 875 447
rect 919 443 923 447
rect 147 431 151 435
rect 487 431 491 435
rect 715 435 719 439
rect 783 435 787 439
rect 827 435 831 439
rect 875 435 879 439
rect 191 423 195 427
rect 555 423 559 427
rect 607 423 611 427
rect 699 427 703 431
rect 791 427 795 431
rect 823 427 827 431
rect 863 427 867 431
rect 791 419 795 423
rect 135 412 139 416
rect 159 412 163 416
rect 183 412 187 416
rect 223 414 227 418
rect 343 414 347 418
rect 447 412 451 416
rect 471 412 475 416
rect 511 414 515 418
rect 615 412 619 416
rect 655 414 659 418
rect 927 412 931 416
rect 111 405 115 409
rect 235 399 239 403
rect 799 401 803 405
rect 959 405 963 409
rect 919 399 923 403
rect 111 387 115 391
rect 175 391 179 395
rect 191 391 195 395
rect 135 378 139 382
rect 147 379 151 383
rect 159 380 163 384
rect 223 388 227 392
rect 343 388 347 392
rect 183 378 187 382
rect 207 383 211 387
rect 427 383 431 387
rect 479 391 483 395
rect 511 388 515 392
rect 607 391 611 395
rect 655 388 659 392
rect 799 388 803 392
rect 935 391 939 395
rect 959 387 963 391
rect 447 380 451 384
rect 459 379 463 383
rect 471 380 475 384
rect 615 380 619 384
rect 627 383 631 387
rect 211 367 215 371
rect 235 367 239 371
rect 243 367 247 371
rect 279 367 283 371
rect 195 355 199 359
rect 331 363 335 367
rect 455 367 459 371
rect 479 367 483 371
rect 487 367 491 371
rect 519 367 523 371
rect 595 367 599 371
rect 687 367 691 371
rect 739 371 743 375
rect 927 380 931 384
rect 323 355 327 359
rect 519 359 523 363
rect 715 363 719 367
rect 647 355 651 359
rect 775 359 779 363
rect 835 359 839 363
rect 207 347 211 351
rect 667 351 671 355
rect 911 351 915 355
rect 215 331 219 335
rect 287 331 291 335
rect 299 331 303 335
rect 323 331 327 335
rect 519 343 523 347
rect 583 343 587 347
rect 687 343 691 347
rect 659 335 663 339
rect 699 335 703 339
rect 775 339 779 343
rect 783 335 787 339
rect 863 343 867 347
rect 831 335 835 339
rect 875 339 879 343
rect 935 343 939 347
rect 903 335 907 339
rect 151 323 155 327
rect 195 323 199 327
rect 207 323 211 327
rect 271 323 275 327
rect 491 323 495 327
rect 547 323 551 327
rect 651 327 655 331
rect 743 327 747 331
rect 667 319 671 323
rect 687 319 691 323
rect 699 319 703 323
rect 863 319 867 323
rect 287 307 291 311
rect 335 307 339 311
rect 743 311 747 315
rect 903 311 907 315
rect 135 300 139 304
rect 159 299 163 303
rect 415 302 419 306
rect 427 299 431 303
rect 439 300 443 304
rect 639 302 643 306
rect 651 303 655 307
rect 767 303 771 307
rect 879 303 883 307
rect 919 307 923 311
rect 927 300 931 304
rect 111 293 115 297
rect 183 292 187 296
rect 311 292 315 296
rect 503 292 507 296
rect 207 283 211 287
rect 423 287 427 291
rect 659 291 663 295
rect 679 292 683 296
rect 807 291 811 295
rect 959 293 963 297
rect 495 287 499 291
rect 863 287 867 291
rect 947 287 951 291
rect 111 275 115 279
rect 311 275 315 279
rect 447 279 451 283
rect 503 279 507 283
rect 679 278 683 282
rect 803 273 807 277
rect 959 275 963 279
rect 135 268 139 272
rect 199 268 203 272
rect 415 268 419 272
rect 439 268 443 272
rect 347 263 351 267
rect 487 267 491 271
rect 639 268 643 272
rect 927 268 931 272
rect 159 255 163 259
rect 175 255 179 259
rect 183 255 187 259
rect 243 251 247 255
rect 295 255 299 259
rect 319 255 323 259
rect 555 259 559 263
rect 647 259 651 263
rect 159 243 163 247
rect 303 247 307 251
rect 463 251 467 255
rect 455 243 456 247
rect 456 243 459 247
rect 487 243 491 247
rect 567 251 571 255
rect 775 255 779 259
rect 935 255 939 259
rect 743 243 747 247
rect 159 235 163 239
rect 243 235 247 239
rect 207 227 211 231
rect 391 231 395 235
rect 239 227 243 231
rect 439 227 443 231
rect 467 231 471 235
rect 567 231 571 235
rect 143 220 147 224
rect 167 220 171 224
rect 191 220 195 224
rect 279 219 283 223
rect 383 220 387 224
rect 407 220 411 224
rect 431 220 435 224
rect 735 220 739 224
rect 775 220 779 224
rect 815 220 819 224
rect 855 220 859 224
rect 903 220 907 224
rect 927 220 931 224
rect 111 213 115 217
rect 475 215 479 219
rect 391 207 395 211
rect 447 207 448 211
rect 448 207 451 211
rect 623 210 627 214
rect 959 213 963 217
rect 111 195 115 199
rect 151 199 155 203
rect 191 199 195 203
rect 143 188 147 192
rect 155 191 159 195
rect 167 188 171 192
rect 179 191 183 195
rect 191 188 195 192
rect 203 187 207 191
rect 303 191 307 195
rect 455 199 459 203
rect 467 199 471 203
rect 535 203 539 207
rect 475 196 479 200
rect 623 196 627 200
rect 743 199 747 203
rect 783 199 787 203
rect 823 199 827 203
rect 887 199 891 203
rect 911 199 915 203
rect 935 199 939 203
rect 959 195 963 199
rect 383 188 387 192
rect 211 183 215 187
rect 395 187 399 191
rect 407 188 411 192
rect 219 183 223 187
rect 431 188 435 192
rect 635 187 639 191
rect 735 188 739 192
rect 747 187 751 191
rect 775 188 779 192
rect 575 179 579 183
rect 599 179 603 183
rect 715 179 719 183
rect 759 179 763 183
rect 815 188 819 192
rect 855 188 859 192
rect 879 187 883 191
rect 903 188 907 192
rect 263 173 267 177
rect 319 167 323 171
rect 335 167 339 171
rect 447 167 451 171
rect 643 167 647 171
rect 747 171 751 175
rect 831 179 835 183
rect 887 179 891 183
rect 927 186 931 190
rect 947 187 951 191
rect 203 159 207 163
rect 271 159 275 163
rect 327 159 331 163
rect 455 151 459 155
rect 487 151 491 155
rect 239 143 243 147
rect 271 143 275 147
rect 211 135 215 139
rect 395 143 399 147
rect 347 131 351 135
rect 423 139 427 143
rect 495 143 499 147
rect 575 151 579 155
rect 687 151 691 155
rect 747 151 751 155
rect 135 124 139 128
rect 111 117 115 121
rect 219 115 223 119
rect 239 124 243 128
rect 367 124 371 128
rect 487 131 491 135
rect 495 124 499 128
rect 623 124 627 128
rect 635 123 639 127
rect 751 124 755 128
rect 959 117 963 121
rect 439 111 443 115
rect 547 111 551 115
rect 759 111 763 115
rect 111 99 115 103
rect 959 99 963 103
rect 135 92 139 96
rect 239 92 243 96
rect 367 92 371 96
rect 495 92 499 96
rect 623 92 627 96
rect 751 92 755 96
<< m3 >>
rect 111 1006 115 1007
rect 111 1001 115 1002
rect 135 1006 139 1007
rect 135 1001 139 1002
rect 319 1006 323 1007
rect 319 1001 323 1002
rect 527 1006 531 1007
rect 527 1001 531 1002
rect 735 1006 739 1007
rect 735 1001 739 1002
rect 927 1006 931 1007
rect 927 1001 931 1002
rect 959 1006 963 1007
rect 959 1001 963 1002
rect 112 994 114 1001
rect 134 1000 140 1001
rect 134 996 135 1000
rect 139 996 140 1000
rect 134 995 140 996
rect 318 1000 324 1001
rect 318 996 319 1000
rect 323 996 324 1000
rect 318 995 324 996
rect 526 1000 532 1001
rect 526 996 527 1000
rect 531 996 532 1000
rect 526 995 532 996
rect 734 1000 740 1001
rect 734 996 735 1000
rect 739 996 740 1000
rect 926 1000 932 1001
rect 926 996 927 1000
rect 931 996 932 1000
rect 734 995 740 996
rect 834 995 840 996
rect 926 995 932 996
rect 110 993 116 994
rect 110 989 111 993
rect 115 989 116 993
rect 834 991 835 995
rect 839 991 840 995
rect 960 994 962 1001
rect 834 990 840 991
rect 958 993 964 994
rect 110 988 116 989
rect 202 979 208 980
rect 110 975 116 976
rect 110 971 111 975
rect 115 971 116 975
rect 202 975 203 979
rect 207 975 208 979
rect 202 974 208 975
rect 110 970 116 971
rect 112 963 114 970
rect 134 968 140 969
rect 134 964 135 968
rect 139 964 140 968
rect 134 963 140 964
rect 111 962 115 963
rect 111 957 115 958
rect 135 962 139 963
rect 135 957 139 958
rect 159 962 163 963
rect 159 957 163 958
rect 183 962 187 963
rect 183 957 187 958
rect 112 914 114 957
rect 136 921 138 957
rect 160 921 162 957
rect 184 921 186 957
rect 134 920 140 921
rect 158 920 164 921
rect 182 920 188 921
rect 134 916 135 920
rect 139 916 140 920
rect 134 915 140 916
rect 146 919 152 920
rect 146 915 147 919
rect 151 915 152 919
rect 158 916 159 920
rect 163 916 164 920
rect 158 915 164 916
rect 170 919 176 920
rect 170 915 171 919
rect 175 915 176 919
rect 182 916 183 920
rect 187 916 188 920
rect 182 915 188 916
rect 146 914 152 915
rect 170 914 178 915
rect 110 913 116 914
rect 110 909 111 913
rect 115 909 116 913
rect 110 908 116 909
rect 110 895 116 896
rect 110 891 111 895
rect 115 891 116 895
rect 110 890 116 891
rect 112 871 114 890
rect 134 888 140 889
rect 134 884 135 888
rect 139 884 140 888
rect 134 883 140 884
rect 126 879 132 880
rect 126 875 127 879
rect 131 875 132 879
rect 126 874 132 875
rect 111 870 115 871
rect 111 865 115 866
rect 112 834 114 865
rect 110 833 116 834
rect 110 829 111 833
rect 115 829 116 833
rect 110 828 116 829
rect 110 815 116 816
rect 110 811 111 815
rect 115 811 116 815
rect 110 810 116 811
rect 112 759 114 810
rect 128 788 130 874
rect 136 871 138 883
rect 135 870 139 871
rect 135 865 139 866
rect 148 864 150 914
rect 172 913 178 914
rect 158 888 164 889
rect 158 884 159 888
rect 163 884 164 888
rect 158 883 164 884
rect 176 883 178 913
rect 190 907 196 908
rect 190 903 191 907
rect 195 903 196 907
rect 190 902 196 903
rect 182 888 188 889
rect 182 884 183 888
rect 187 884 188 888
rect 182 883 188 884
rect 160 871 162 883
rect 168 881 178 883
rect 159 870 163 871
rect 159 865 163 866
rect 146 863 152 864
rect 146 859 147 863
rect 151 859 152 863
rect 146 858 152 859
rect 150 855 156 856
rect 150 851 151 855
rect 155 851 156 855
rect 150 850 156 851
rect 126 787 132 788
rect 126 783 127 787
rect 131 783 132 787
rect 126 782 132 783
rect 111 758 115 759
rect 111 753 115 754
rect 135 758 139 759
rect 135 753 139 754
rect 112 710 114 753
rect 136 717 138 753
rect 134 716 140 717
rect 134 712 135 716
rect 139 712 140 716
rect 134 711 140 712
rect 110 709 116 710
rect 110 705 111 709
rect 115 705 116 709
rect 110 704 116 705
rect 142 703 148 704
rect 142 699 143 703
rect 147 699 148 703
rect 142 698 148 699
rect 110 691 116 692
rect 110 687 111 691
rect 115 687 116 691
rect 110 686 116 687
rect 112 659 114 686
rect 134 684 140 685
rect 134 680 135 684
rect 139 680 140 684
rect 134 679 140 680
rect 136 659 138 679
rect 144 668 146 698
rect 152 676 154 850
rect 168 848 170 881
rect 184 871 186 883
rect 192 880 194 902
rect 190 879 196 880
rect 190 875 191 879
rect 195 875 196 879
rect 190 874 196 875
rect 175 870 179 871
rect 175 865 179 866
rect 183 870 187 871
rect 183 865 187 866
rect 166 847 172 848
rect 166 843 167 847
rect 171 843 172 847
rect 166 842 172 843
rect 176 841 178 865
rect 174 840 180 841
rect 174 836 175 840
rect 179 836 180 840
rect 174 835 180 836
rect 158 816 164 817
rect 158 812 159 816
rect 163 812 164 816
rect 158 811 164 812
rect 160 759 162 811
rect 204 808 206 974
rect 318 968 324 969
rect 318 964 319 968
rect 323 964 324 968
rect 318 963 324 964
rect 526 968 532 969
rect 526 964 527 968
rect 531 964 532 968
rect 526 963 532 964
rect 734 968 740 969
rect 734 964 735 968
rect 739 964 740 968
rect 734 963 740 964
rect 758 967 764 968
rect 758 963 759 967
rect 763 963 764 967
rect 231 962 235 963
rect 231 957 235 958
rect 311 962 315 963
rect 311 957 315 958
rect 319 962 323 963
rect 455 962 459 963
rect 319 957 323 958
rect 426 959 432 960
rect 232 921 234 957
rect 286 951 292 952
rect 286 947 287 951
rect 291 950 292 951
rect 298 951 304 952
rect 291 947 294 950
rect 286 946 294 947
rect 298 947 299 951
rect 303 947 304 951
rect 298 946 304 947
rect 230 920 236 921
rect 222 919 228 920
rect 222 915 223 919
rect 227 915 228 919
rect 230 916 231 920
rect 235 916 236 920
rect 230 915 236 916
rect 250 919 256 920
rect 250 915 251 919
rect 255 915 256 919
rect 222 914 228 915
rect 250 914 256 915
rect 224 856 226 914
rect 238 907 244 908
rect 238 903 239 907
rect 243 903 244 907
rect 238 902 244 903
rect 230 888 236 889
rect 230 884 231 888
rect 235 884 236 888
rect 230 883 236 884
rect 232 871 234 883
rect 231 870 235 871
rect 231 865 235 866
rect 222 855 228 856
rect 222 851 223 855
rect 227 851 228 855
rect 222 850 228 851
rect 230 855 236 856
rect 230 851 231 855
rect 235 851 236 855
rect 230 850 236 851
rect 202 807 208 808
rect 202 803 203 807
rect 207 803 208 807
rect 202 802 208 803
rect 198 779 204 780
rect 198 775 199 779
rect 203 775 204 779
rect 198 774 204 775
rect 159 758 163 759
rect 159 753 163 754
rect 175 758 179 759
rect 175 753 179 754
rect 176 709 178 753
rect 200 732 202 774
rect 232 732 234 850
rect 240 756 242 902
rect 252 900 254 914
rect 250 899 256 900
rect 250 895 251 899
rect 255 895 256 899
rect 250 894 256 895
rect 274 879 280 880
rect 274 875 275 879
rect 279 875 280 879
rect 274 874 280 875
rect 276 828 278 874
rect 274 827 280 828
rect 274 823 275 827
rect 279 823 280 827
rect 274 822 280 823
rect 276 796 278 822
rect 274 795 280 796
rect 274 791 275 795
rect 279 791 280 795
rect 274 790 280 791
rect 292 771 294 946
rect 300 928 302 946
rect 298 927 304 928
rect 298 923 299 927
rect 303 923 304 927
rect 298 922 304 923
rect 298 919 304 920
rect 298 915 299 919
rect 303 915 304 919
rect 298 914 304 915
rect 300 780 302 914
rect 312 913 314 957
rect 426 955 427 959
rect 431 955 432 959
rect 455 957 459 958
rect 519 962 523 963
rect 519 957 523 958
rect 527 962 531 963
rect 527 957 531 958
rect 583 962 587 963
rect 583 957 587 958
rect 647 962 651 963
rect 647 957 651 958
rect 711 962 715 963
rect 711 957 715 958
rect 735 962 739 963
rect 758 962 764 963
rect 767 962 771 963
rect 735 957 739 958
rect 426 954 432 955
rect 318 951 324 952
rect 318 947 319 951
rect 323 947 324 951
rect 318 946 324 947
rect 310 912 316 913
rect 310 908 311 912
rect 315 908 316 912
rect 310 907 316 908
rect 310 895 316 896
rect 310 891 311 895
rect 315 891 316 895
rect 310 890 316 891
rect 312 871 314 890
rect 311 870 315 871
rect 311 865 315 866
rect 310 793 316 794
rect 310 789 311 793
rect 315 789 316 793
rect 310 788 316 789
rect 298 779 304 780
rect 298 775 299 779
rect 303 775 304 779
rect 298 774 304 775
rect 292 769 298 771
rect 279 758 283 759
rect 238 755 244 756
rect 238 751 239 755
rect 243 751 244 755
rect 279 753 283 754
rect 238 750 244 751
rect 198 731 204 732
rect 198 727 199 731
rect 203 727 204 731
rect 198 726 204 727
rect 230 731 236 732
rect 230 727 231 731
rect 235 727 236 731
rect 230 726 236 727
rect 174 708 180 709
rect 174 704 175 708
rect 179 704 180 708
rect 174 703 180 704
rect 174 682 180 683
rect 174 678 175 682
rect 179 678 180 682
rect 174 677 180 678
rect 150 675 156 676
rect 150 671 151 675
rect 155 671 156 675
rect 150 670 156 671
rect 142 667 148 668
rect 142 663 143 667
rect 147 663 148 667
rect 142 662 148 663
rect 111 658 115 659
rect 111 653 115 654
rect 135 658 139 659
rect 135 653 139 654
rect 112 622 114 653
rect 110 621 116 622
rect 110 617 111 621
rect 115 617 116 621
rect 110 616 116 617
rect 110 603 116 604
rect 110 599 111 603
rect 115 599 116 603
rect 110 598 116 599
rect 112 547 114 598
rect 144 564 146 662
rect 176 659 178 677
rect 159 658 163 659
rect 159 653 163 654
rect 175 658 179 659
rect 175 653 179 654
rect 160 622 162 653
rect 158 621 164 622
rect 158 617 159 621
rect 163 617 164 621
rect 158 616 164 617
rect 158 604 164 605
rect 158 600 159 604
rect 163 600 164 604
rect 158 599 164 600
rect 134 563 140 564
rect 134 559 135 563
rect 139 559 140 563
rect 134 558 140 559
rect 144 563 152 564
rect 144 559 147 563
rect 151 559 152 563
rect 144 558 152 559
rect 111 546 115 547
rect 111 541 115 542
rect 112 490 114 541
rect 136 512 138 558
rect 144 520 146 558
rect 160 547 162 599
rect 200 592 202 726
rect 280 717 282 753
rect 296 740 298 769
rect 312 759 314 788
rect 320 764 322 946
rect 370 911 376 912
rect 370 907 371 911
rect 375 907 376 911
rect 370 906 376 907
rect 338 875 344 876
rect 338 871 339 875
rect 343 871 344 875
rect 327 870 331 871
rect 338 870 344 871
rect 346 875 352 876
rect 346 871 347 875
rect 351 871 352 875
rect 346 870 352 871
rect 327 865 331 866
rect 328 840 330 865
rect 340 860 342 870
rect 338 859 344 860
rect 338 855 339 859
rect 343 855 344 859
rect 338 854 344 855
rect 326 839 332 840
rect 326 835 327 839
rect 331 835 332 839
rect 326 834 332 835
rect 348 828 350 870
rect 358 847 364 848
rect 358 843 359 847
rect 363 843 364 847
rect 358 842 364 843
rect 346 827 352 828
rect 346 823 347 827
rect 351 823 352 827
rect 346 822 352 823
rect 318 763 324 764
rect 318 759 319 763
rect 323 759 324 763
rect 303 758 307 759
rect 303 753 307 754
rect 311 758 315 759
rect 318 758 324 759
rect 327 758 331 759
rect 311 753 315 754
rect 327 753 331 754
rect 351 758 355 759
rect 351 753 355 754
rect 294 739 300 740
rect 294 735 295 739
rect 299 735 300 739
rect 294 734 300 735
rect 304 717 306 753
rect 314 723 320 724
rect 314 719 315 723
rect 319 719 320 723
rect 314 718 320 719
rect 278 716 284 717
rect 302 716 308 717
rect 278 712 279 716
rect 283 712 284 716
rect 278 711 284 712
rect 290 715 296 716
rect 290 711 291 715
rect 295 714 296 715
rect 295 711 298 714
rect 302 712 303 716
rect 307 712 308 716
rect 316 715 318 718
rect 328 717 330 753
rect 352 719 354 753
rect 360 748 362 842
rect 372 795 374 906
rect 378 903 384 904
rect 378 899 379 903
rect 383 899 384 903
rect 378 898 384 899
rect 380 852 382 898
rect 428 884 430 954
rect 442 951 448 952
rect 442 947 443 951
rect 447 947 448 951
rect 442 946 448 947
rect 426 883 432 884
rect 426 879 427 883
rect 431 879 432 883
rect 426 878 432 879
rect 434 879 440 880
rect 434 875 435 879
rect 439 875 440 879
rect 432 874 440 875
rect 432 873 438 874
rect 378 851 384 852
rect 378 847 379 851
rect 383 847 384 851
rect 378 846 384 847
rect 386 851 392 852
rect 386 847 387 851
rect 391 847 392 851
rect 386 846 392 847
rect 388 843 390 846
rect 384 841 390 843
rect 384 804 386 841
rect 382 803 388 804
rect 382 799 383 803
rect 387 799 388 803
rect 382 798 388 799
rect 368 793 374 795
rect 368 788 370 793
rect 366 787 372 788
rect 366 783 367 787
rect 371 783 372 787
rect 366 782 372 783
rect 374 787 380 788
rect 374 783 375 787
rect 379 783 380 787
rect 374 782 380 783
rect 366 779 372 780
rect 366 775 367 779
rect 371 775 372 779
rect 366 774 372 775
rect 368 764 370 774
rect 366 763 372 764
rect 366 759 367 763
rect 371 759 372 763
rect 366 758 372 759
rect 358 747 364 748
rect 358 743 359 747
rect 363 743 364 747
rect 358 742 364 743
rect 376 740 378 782
rect 432 772 434 873
rect 444 788 446 946
rect 456 921 458 957
rect 520 921 522 957
rect 584 921 586 957
rect 648 921 650 957
rect 712 921 714 957
rect 454 920 460 921
rect 518 920 524 921
rect 582 920 588 921
rect 646 920 652 921
rect 710 920 716 921
rect 454 916 455 920
rect 459 916 460 920
rect 454 915 460 916
rect 466 919 472 920
rect 466 915 467 919
rect 471 918 472 919
rect 471 915 474 918
rect 518 916 519 920
rect 523 916 524 920
rect 518 915 524 916
rect 530 919 536 920
rect 530 915 531 919
rect 535 915 536 919
rect 582 916 583 920
rect 587 916 588 920
rect 582 915 588 916
rect 630 919 636 920
rect 630 915 631 919
rect 635 915 636 919
rect 646 916 647 920
rect 651 916 652 920
rect 646 915 652 916
rect 666 919 672 920
rect 666 915 667 919
rect 671 915 672 919
rect 710 916 711 920
rect 715 916 716 920
rect 710 915 716 916
rect 722 919 728 920
rect 722 915 723 919
rect 727 918 728 919
rect 727 915 730 918
rect 466 914 474 915
rect 530 914 536 915
rect 630 914 636 915
rect 666 914 672 915
rect 722 914 730 915
rect 458 888 464 889
rect 458 884 459 888
rect 463 884 464 888
rect 458 883 464 884
rect 460 871 462 883
rect 451 870 455 871
rect 451 865 455 866
rect 459 870 463 871
rect 459 865 463 866
rect 452 836 454 865
rect 450 835 456 836
rect 450 831 451 835
rect 455 831 456 835
rect 450 830 456 831
rect 450 816 456 817
rect 450 812 451 816
rect 455 812 456 816
rect 450 811 456 812
rect 442 787 448 788
rect 442 783 443 787
rect 447 783 448 787
rect 442 782 448 783
rect 430 771 436 772
rect 430 767 431 771
rect 435 767 436 771
rect 444 768 446 782
rect 430 766 436 767
rect 442 767 448 768
rect 442 763 443 767
rect 447 763 448 767
rect 442 762 448 763
rect 452 759 454 811
rect 472 808 474 914
rect 510 903 516 904
rect 510 899 511 903
rect 515 899 516 903
rect 510 898 516 899
rect 470 807 476 808
rect 470 803 471 807
rect 475 803 476 807
rect 470 802 476 803
rect 486 787 492 788
rect 486 783 487 787
rect 491 783 492 787
rect 486 782 492 783
rect 383 758 387 759
rect 383 753 387 754
rect 415 758 419 759
rect 415 753 419 754
rect 439 758 443 759
rect 439 753 443 754
rect 451 758 455 759
rect 451 753 455 754
rect 463 758 467 759
rect 463 753 467 754
rect 374 739 380 740
rect 374 735 375 739
rect 379 735 380 739
rect 374 734 380 735
rect 376 720 378 734
rect 374 719 380 720
rect 350 718 356 719
rect 326 716 332 717
rect 316 713 322 715
rect 302 711 308 712
rect 290 710 298 711
rect 286 703 292 704
rect 286 699 287 703
rect 291 699 292 703
rect 286 698 292 699
rect 278 684 284 685
rect 278 680 279 684
rect 283 680 284 684
rect 278 679 284 680
rect 280 659 282 679
rect 279 658 283 659
rect 279 653 283 654
rect 274 643 280 644
rect 274 639 275 643
rect 279 639 280 643
rect 274 638 280 639
rect 262 631 268 632
rect 262 627 263 631
rect 267 627 268 631
rect 262 626 268 627
rect 230 611 236 612
rect 230 607 231 611
rect 235 607 236 611
rect 230 606 236 607
rect 198 591 204 592
rect 198 587 199 591
rect 203 587 204 591
rect 198 586 204 587
rect 151 546 155 547
rect 151 541 155 542
rect 159 546 163 547
rect 159 541 163 542
rect 142 519 148 520
rect 142 515 143 519
rect 147 515 148 519
rect 142 514 148 515
rect 136 511 144 512
rect 136 507 139 511
rect 143 507 144 511
rect 136 506 144 507
rect 136 505 142 506
rect 110 489 116 490
rect 110 485 111 489
rect 115 485 116 489
rect 110 484 116 485
rect 140 475 142 505
rect 152 489 154 541
rect 174 495 180 496
rect 174 491 175 495
rect 179 491 180 495
rect 174 490 180 491
rect 150 488 156 489
rect 150 484 151 488
rect 155 484 156 488
rect 150 483 156 484
rect 140 473 146 475
rect 110 471 116 472
rect 110 467 111 471
rect 115 467 116 471
rect 110 466 116 467
rect 112 447 114 466
rect 111 446 115 447
rect 111 441 115 442
rect 135 446 139 447
rect 135 441 139 442
rect 112 410 114 441
rect 136 417 138 441
rect 144 436 146 473
rect 150 462 156 463
rect 150 458 151 462
rect 155 458 156 462
rect 150 457 156 458
rect 152 447 154 457
rect 151 446 155 447
rect 151 441 155 442
rect 159 446 163 447
rect 159 441 163 442
rect 144 435 152 436
rect 144 433 147 435
rect 146 431 147 433
rect 151 431 152 435
rect 146 430 152 431
rect 134 416 140 417
rect 134 412 135 416
rect 139 412 140 416
rect 134 411 140 412
rect 110 409 116 410
rect 110 405 111 409
rect 115 405 116 409
rect 110 404 116 405
rect 110 391 116 392
rect 110 387 111 391
rect 115 387 116 391
rect 110 386 116 387
rect 112 355 114 386
rect 148 384 150 430
rect 160 417 162 441
rect 158 416 164 417
rect 158 412 159 416
rect 163 412 164 416
rect 158 411 164 412
rect 176 396 178 490
rect 232 452 234 606
rect 238 563 244 564
rect 238 559 239 563
rect 243 559 244 563
rect 264 563 266 626
rect 276 613 278 638
rect 275 612 279 613
rect 274 607 275 612
rect 279 607 280 612
rect 288 611 290 698
rect 296 652 298 710
rect 302 684 308 685
rect 302 680 303 684
rect 307 680 308 684
rect 302 679 308 680
rect 304 659 306 679
rect 320 668 322 713
rect 326 712 327 716
rect 331 712 332 716
rect 326 711 332 712
rect 338 715 344 716
rect 338 711 339 715
rect 343 714 344 715
rect 350 714 351 718
rect 355 714 356 718
rect 374 715 375 719
rect 379 715 380 719
rect 384 717 386 753
rect 416 719 418 753
rect 414 718 420 719
rect 374 714 380 715
rect 382 716 388 717
rect 343 711 346 714
rect 350 713 356 714
rect 382 712 383 716
rect 387 712 388 716
rect 382 711 388 712
rect 406 715 412 716
rect 406 711 407 715
rect 411 711 412 715
rect 414 714 415 718
rect 419 714 420 718
rect 440 717 442 753
rect 450 747 456 748
rect 450 743 451 747
rect 455 743 456 747
rect 450 742 456 743
rect 414 713 420 714
rect 438 716 444 717
rect 452 716 454 742
rect 464 717 466 753
rect 478 747 484 748
rect 478 743 479 747
rect 483 743 484 747
rect 478 742 484 743
rect 462 716 468 717
rect 438 712 439 716
rect 443 712 444 716
rect 438 711 444 712
rect 450 715 456 716
rect 450 711 451 715
rect 455 711 456 715
rect 462 712 463 716
rect 467 712 468 716
rect 462 711 468 712
rect 338 710 346 711
rect 406 710 412 711
rect 450 710 456 711
rect 326 684 332 685
rect 326 680 327 684
rect 331 680 332 684
rect 326 679 332 680
rect 318 667 324 668
rect 318 663 319 667
rect 323 663 324 667
rect 318 662 324 663
rect 328 659 330 679
rect 303 658 307 659
rect 303 653 307 654
rect 327 658 331 659
rect 327 653 331 654
rect 294 651 300 652
rect 294 647 295 651
rect 299 647 300 651
rect 294 646 300 647
rect 304 629 306 653
rect 344 650 346 710
rect 358 703 364 704
rect 358 699 359 703
rect 363 699 364 703
rect 358 698 364 699
rect 390 703 396 704
rect 390 699 391 703
rect 395 699 396 703
rect 390 698 396 699
rect 350 684 356 685
rect 350 680 351 684
rect 355 680 356 684
rect 350 679 356 680
rect 352 659 354 679
rect 360 676 362 698
rect 382 684 388 685
rect 382 680 383 684
rect 387 680 388 684
rect 382 679 388 680
rect 358 675 364 676
rect 358 671 359 675
rect 363 671 364 675
rect 358 670 364 671
rect 384 659 386 679
rect 351 658 355 659
rect 351 653 355 654
rect 383 658 387 659
rect 383 653 387 654
rect 336 648 346 650
rect 336 636 338 648
rect 334 635 340 636
rect 334 631 335 635
rect 339 631 340 635
rect 334 630 340 631
rect 302 628 308 629
rect 302 624 303 628
rect 307 624 308 628
rect 302 623 308 624
rect 358 611 364 612
rect 288 609 298 611
rect 274 606 280 607
rect 276 603 278 606
rect 286 604 292 605
rect 286 600 287 604
rect 291 600 292 604
rect 286 599 292 600
rect 278 591 284 592
rect 278 587 279 591
rect 283 587 284 591
rect 278 586 284 587
rect 280 572 282 586
rect 278 571 284 572
rect 278 567 279 571
rect 283 567 284 571
rect 278 566 284 567
rect 264 561 270 563
rect 238 558 244 559
rect 240 544 242 558
rect 255 546 259 547
rect 238 543 244 544
rect 238 539 239 543
rect 243 539 244 543
rect 255 541 259 542
rect 238 538 244 539
rect 256 497 258 541
rect 254 496 260 497
rect 268 496 270 561
rect 288 547 290 599
rect 296 576 298 609
rect 358 607 359 611
rect 363 607 364 611
rect 358 606 364 607
rect 326 595 332 596
rect 326 594 327 595
rect 320 592 327 594
rect 294 575 300 576
rect 294 571 295 575
rect 299 571 300 575
rect 294 570 300 571
rect 279 546 283 547
rect 279 541 283 542
rect 287 546 291 547
rect 287 541 291 542
rect 303 546 307 547
rect 303 541 307 542
rect 280 497 282 541
rect 304 497 306 541
rect 310 503 316 504
rect 310 499 311 503
rect 315 499 316 503
rect 310 498 316 499
rect 278 496 284 497
rect 302 496 308 497
rect 254 492 255 496
rect 259 492 260 496
rect 254 491 260 492
rect 266 495 272 496
rect 266 491 267 495
rect 271 491 272 495
rect 278 492 279 496
rect 283 492 284 496
rect 278 491 284 492
rect 290 495 296 496
rect 290 491 291 495
rect 295 491 296 495
rect 302 492 303 496
rect 307 492 308 496
rect 302 491 308 492
rect 266 490 272 491
rect 288 490 296 491
rect 288 489 294 490
rect 288 486 290 489
rect 312 486 314 498
rect 320 488 322 592
rect 326 591 327 592
rect 331 591 332 595
rect 326 590 332 591
rect 350 575 356 576
rect 350 571 351 575
rect 355 571 356 575
rect 350 570 356 571
rect 327 546 331 547
rect 327 541 331 542
rect 328 497 330 541
rect 326 496 332 497
rect 326 492 327 496
rect 331 492 332 496
rect 326 491 332 492
rect 352 488 354 570
rect 360 536 362 606
rect 382 583 388 584
rect 382 579 383 583
rect 387 579 388 583
rect 382 578 388 579
rect 384 564 386 578
rect 382 563 388 564
rect 382 559 383 563
rect 387 559 388 563
rect 382 558 388 559
rect 379 546 383 547
rect 379 541 383 542
rect 370 539 376 540
rect 358 535 364 536
rect 358 531 359 535
rect 363 531 364 535
rect 370 535 371 539
rect 375 535 376 539
rect 370 534 376 535
rect 358 530 364 531
rect 372 512 374 534
rect 370 511 376 512
rect 370 507 371 511
rect 375 507 376 511
rect 370 506 376 507
rect 380 489 382 541
rect 392 540 394 698
rect 408 696 410 710
rect 422 703 428 704
rect 422 699 423 703
rect 427 699 428 703
rect 422 698 428 699
rect 446 703 452 704
rect 446 699 447 703
rect 451 699 452 703
rect 446 698 452 699
rect 406 695 412 696
rect 406 691 407 695
rect 411 691 412 695
rect 406 690 412 691
rect 408 651 410 690
rect 414 684 420 685
rect 414 680 415 684
rect 419 680 420 684
rect 414 679 420 680
rect 416 659 418 679
rect 415 658 419 659
rect 415 653 419 654
rect 408 649 414 651
rect 412 568 414 649
rect 410 567 416 568
rect 410 563 411 567
rect 415 563 416 567
rect 410 562 416 563
rect 390 539 396 540
rect 390 535 391 539
rect 395 535 396 539
rect 390 534 396 535
rect 424 512 426 698
rect 438 684 444 685
rect 438 680 439 684
rect 443 680 444 684
rect 438 679 444 680
rect 440 659 442 679
rect 439 658 443 659
rect 439 653 443 654
rect 430 635 436 636
rect 430 631 431 635
rect 435 631 436 635
rect 430 630 436 631
rect 422 511 428 512
rect 422 507 423 511
rect 427 507 428 511
rect 422 506 428 507
rect 378 488 384 489
rect 432 488 434 630
rect 438 581 444 582
rect 438 577 439 581
rect 443 577 444 581
rect 438 576 444 577
rect 440 547 442 576
rect 439 546 443 547
rect 439 541 443 542
rect 438 531 444 532
rect 438 527 439 531
rect 443 527 444 531
rect 438 526 444 527
rect 280 484 290 486
rect 304 484 314 486
rect 318 487 324 488
rect 278 483 284 484
rect 278 479 279 483
rect 283 479 284 483
rect 278 478 284 479
rect 302 483 308 484
rect 302 479 303 483
rect 307 479 308 483
rect 318 483 319 487
rect 323 483 324 487
rect 318 482 324 483
rect 350 487 356 488
rect 350 483 351 487
rect 355 483 356 487
rect 378 484 379 488
rect 383 484 384 488
rect 378 483 384 484
rect 430 487 436 488
rect 430 483 431 487
rect 435 483 436 487
rect 350 482 356 483
rect 430 482 436 483
rect 302 478 308 479
rect 378 469 384 470
rect 378 465 379 469
rect 383 465 384 469
rect 254 464 260 465
rect 254 460 255 464
rect 259 460 260 464
rect 254 459 260 460
rect 278 464 284 465
rect 278 460 279 464
rect 283 460 284 464
rect 278 459 284 460
rect 302 464 308 465
rect 302 460 303 464
rect 307 460 308 464
rect 302 459 308 460
rect 326 464 332 465
rect 378 464 384 465
rect 326 460 327 464
rect 331 460 332 464
rect 326 459 332 460
rect 230 451 236 452
rect 230 447 231 451
rect 235 447 236 451
rect 256 447 258 459
rect 280 447 282 459
rect 304 447 306 459
rect 328 447 330 459
rect 380 447 382 464
rect 440 456 442 526
rect 448 480 450 698
rect 462 684 468 685
rect 462 680 463 684
rect 467 680 468 684
rect 462 679 468 680
rect 464 659 466 679
rect 455 658 459 659
rect 455 653 459 654
rect 463 658 467 659
rect 463 653 467 654
rect 456 628 458 653
rect 466 647 472 648
rect 466 643 467 647
rect 471 643 472 647
rect 466 642 472 643
rect 454 627 460 628
rect 454 623 455 627
rect 459 623 460 627
rect 454 622 460 623
rect 454 567 460 568
rect 454 563 455 567
rect 459 563 460 567
rect 454 562 460 563
rect 456 552 458 562
rect 454 551 460 552
rect 454 547 455 551
rect 459 547 460 551
rect 454 546 460 547
rect 468 532 470 642
rect 480 600 482 742
rect 488 708 490 782
rect 512 764 514 898
rect 532 896 534 914
rect 538 907 544 908
rect 538 903 539 907
rect 543 903 544 907
rect 538 902 544 903
rect 530 895 536 896
rect 530 891 531 895
rect 535 891 536 895
rect 530 890 536 891
rect 518 888 524 889
rect 518 884 519 888
rect 523 884 524 888
rect 518 883 524 884
rect 520 871 522 883
rect 519 870 523 871
rect 519 865 523 866
rect 540 864 542 902
rect 582 888 588 889
rect 582 884 583 888
rect 587 884 588 888
rect 582 883 588 884
rect 584 871 586 883
rect 575 870 579 871
rect 575 865 579 866
rect 583 870 587 871
rect 583 865 587 866
rect 538 863 544 864
rect 538 859 539 863
rect 543 859 544 863
rect 538 858 544 859
rect 526 855 532 856
rect 518 851 524 852
rect 518 847 519 851
rect 523 847 524 851
rect 526 851 527 855
rect 531 851 532 855
rect 526 850 532 851
rect 518 846 524 847
rect 520 832 522 846
rect 518 831 524 832
rect 518 827 519 831
rect 523 827 524 831
rect 518 826 524 827
rect 528 772 530 850
rect 540 772 542 858
rect 562 847 568 848
rect 562 843 563 847
rect 567 843 568 847
rect 562 842 568 843
rect 554 799 560 800
rect 554 795 555 799
rect 559 795 560 799
rect 554 794 560 795
rect 556 772 558 794
rect 526 771 532 772
rect 526 767 527 771
rect 531 767 532 771
rect 526 766 532 767
rect 538 771 544 772
rect 538 767 539 771
rect 543 767 544 771
rect 538 766 544 767
rect 554 771 560 772
rect 554 767 555 771
rect 559 767 560 771
rect 554 766 560 767
rect 510 763 516 764
rect 510 759 511 763
rect 515 759 516 763
rect 495 758 499 759
rect 510 758 516 759
rect 495 753 499 754
rect 512 755 514 758
rect 528 756 530 766
rect 543 758 547 759
rect 526 755 532 756
rect 512 753 518 755
rect 496 719 498 753
rect 506 743 512 744
rect 506 739 507 743
rect 511 739 512 743
rect 506 738 512 739
rect 508 720 510 738
rect 516 736 518 753
rect 526 751 527 755
rect 531 751 532 755
rect 543 753 547 754
rect 550 755 556 756
rect 526 750 532 751
rect 514 735 520 736
rect 514 731 515 735
rect 519 731 520 735
rect 514 730 520 731
rect 506 719 512 720
rect 494 718 500 719
rect 494 714 495 718
rect 499 714 500 718
rect 506 715 507 719
rect 511 715 512 719
rect 506 714 512 715
rect 494 713 500 714
rect 544 709 546 753
rect 550 751 551 755
rect 555 751 556 755
rect 550 750 556 751
rect 552 736 554 750
rect 564 736 566 842
rect 576 841 578 865
rect 574 840 580 841
rect 574 836 575 840
rect 579 836 580 840
rect 574 835 580 836
rect 586 827 592 828
rect 586 823 587 827
rect 591 823 592 827
rect 586 822 592 823
rect 588 812 590 822
rect 594 819 600 820
rect 594 815 595 819
rect 599 815 600 819
rect 594 814 600 815
rect 586 811 592 812
rect 574 808 580 809
rect 574 804 575 808
rect 579 804 580 808
rect 586 807 587 811
rect 591 807 592 811
rect 586 806 592 807
rect 574 803 580 804
rect 576 759 578 803
rect 588 797 590 806
rect 587 796 591 797
rect 587 791 591 792
rect 575 758 579 759
rect 575 753 579 754
rect 596 740 598 814
rect 632 812 634 914
rect 654 907 660 908
rect 654 903 655 907
rect 659 903 660 907
rect 654 902 660 903
rect 646 888 652 889
rect 646 884 647 888
rect 651 884 652 888
rect 646 883 652 884
rect 648 871 650 883
rect 639 870 643 871
rect 639 865 643 866
rect 647 870 651 871
rect 647 865 651 866
rect 640 830 642 865
rect 656 856 658 902
rect 654 855 660 856
rect 654 851 655 855
rect 659 851 660 855
rect 654 850 660 851
rect 638 829 644 830
rect 638 825 639 829
rect 643 825 644 829
rect 638 824 644 825
rect 638 816 644 817
rect 638 812 639 816
rect 643 812 644 816
rect 630 811 636 812
rect 638 811 644 812
rect 630 807 631 811
rect 635 807 636 811
rect 630 806 636 807
rect 626 783 632 784
rect 626 779 627 783
rect 631 779 632 783
rect 626 778 632 779
rect 628 764 630 778
rect 626 763 632 764
rect 626 759 627 763
rect 631 759 632 763
rect 640 759 642 811
rect 626 758 632 759
rect 639 758 643 759
rect 639 753 643 754
rect 655 758 659 759
rect 668 756 670 914
rect 702 907 708 908
rect 702 903 703 907
rect 707 903 708 907
rect 702 902 708 903
rect 704 880 706 902
rect 710 888 716 889
rect 710 884 711 888
rect 715 884 716 888
rect 710 883 716 884
rect 702 879 708 880
rect 702 875 703 879
rect 707 875 708 879
rect 702 874 708 875
rect 704 856 706 874
rect 712 871 714 883
rect 728 872 730 914
rect 726 871 732 872
rect 711 870 715 871
rect 726 867 727 871
rect 731 867 732 871
rect 726 866 732 867
rect 711 865 715 866
rect 728 860 730 866
rect 726 859 732 860
rect 702 855 708 856
rect 702 851 703 855
rect 707 851 708 855
rect 726 855 727 859
rect 731 855 732 859
rect 726 854 732 855
rect 702 850 708 851
rect 738 799 744 800
rect 738 795 739 799
rect 743 795 744 799
rect 738 794 744 795
rect 682 771 688 772
rect 682 767 683 771
rect 687 767 688 771
rect 682 766 688 767
rect 655 753 659 754
rect 666 755 672 756
rect 594 739 600 740
rect 550 735 556 736
rect 550 731 551 735
rect 555 731 556 735
rect 550 730 556 731
rect 562 735 568 736
rect 562 731 563 735
rect 567 731 568 735
rect 594 735 595 739
rect 599 735 600 739
rect 594 734 600 735
rect 562 730 568 731
rect 542 708 548 709
rect 486 707 492 708
rect 486 703 487 707
rect 491 703 492 707
rect 542 704 543 708
rect 547 704 548 708
rect 542 703 548 704
rect 486 702 492 703
rect 486 699 492 700
rect 486 695 487 699
rect 491 695 492 699
rect 486 694 492 695
rect 542 694 548 695
rect 478 599 484 600
rect 478 595 479 599
rect 483 595 484 599
rect 478 594 484 595
rect 488 560 490 694
rect 542 690 543 694
rect 547 690 548 694
rect 542 689 548 690
rect 494 684 500 685
rect 494 680 495 684
rect 499 680 500 684
rect 494 679 500 680
rect 496 659 498 679
rect 544 659 546 689
rect 564 676 566 730
rect 656 717 658 753
rect 666 751 667 755
rect 671 751 672 755
rect 666 750 672 751
rect 684 740 686 766
rect 695 758 699 759
rect 695 753 699 754
rect 710 755 716 756
rect 682 739 688 740
rect 682 735 683 739
rect 687 735 688 739
rect 682 734 688 735
rect 654 716 660 717
rect 654 712 655 716
rect 659 712 660 716
rect 654 711 660 712
rect 696 709 698 753
rect 710 751 711 755
rect 715 751 716 755
rect 710 750 716 751
rect 712 732 714 750
rect 710 731 716 732
rect 710 727 711 731
rect 715 727 716 731
rect 710 726 716 727
rect 694 708 700 709
rect 694 704 695 708
rect 699 704 700 708
rect 662 703 668 704
rect 694 703 700 704
rect 662 699 663 703
rect 667 699 668 703
rect 662 698 668 699
rect 654 684 660 685
rect 654 680 655 684
rect 659 680 660 684
rect 654 679 660 680
rect 562 675 568 676
rect 562 671 563 675
rect 567 671 568 675
rect 562 670 568 671
rect 656 659 658 679
rect 664 660 666 698
rect 694 682 700 683
rect 694 678 695 682
rect 699 678 700 682
rect 694 677 700 678
rect 670 667 676 668
rect 670 663 671 667
rect 675 663 676 667
rect 670 662 676 663
rect 662 659 668 660
rect 495 658 499 659
rect 495 653 499 654
rect 543 658 547 659
rect 543 653 547 654
rect 559 658 563 659
rect 559 653 563 654
rect 583 658 587 659
rect 583 653 587 654
rect 647 658 651 659
rect 647 653 651 654
rect 655 658 659 659
rect 662 655 663 659
rect 667 655 668 659
rect 662 654 668 655
rect 655 653 659 654
rect 560 629 562 653
rect 566 639 572 640
rect 566 635 567 639
rect 571 635 572 639
rect 566 634 572 635
rect 558 628 564 629
rect 558 624 559 628
rect 563 624 564 628
rect 558 623 564 624
rect 510 615 516 616
rect 510 611 511 615
rect 515 614 516 615
rect 538 615 544 616
rect 538 614 539 615
rect 515 612 539 614
rect 515 611 516 612
rect 510 610 516 611
rect 538 611 539 612
rect 543 611 544 615
rect 538 610 544 611
rect 568 608 570 634
rect 584 629 586 653
rect 594 651 600 652
rect 594 647 595 651
rect 599 647 600 651
rect 594 646 600 647
rect 638 651 644 652
rect 638 647 639 651
rect 643 647 644 651
rect 638 646 644 647
rect 582 628 588 629
rect 582 624 583 628
rect 587 624 588 628
rect 582 623 588 624
rect 550 607 556 608
rect 550 603 551 607
rect 555 603 556 607
rect 550 602 556 603
rect 566 607 572 608
rect 566 603 567 607
rect 571 603 572 607
rect 566 602 572 603
rect 552 564 554 602
rect 558 596 564 597
rect 582 596 588 597
rect 596 596 598 646
rect 618 643 624 644
rect 618 639 619 643
rect 623 639 624 643
rect 618 638 624 639
rect 606 635 612 636
rect 606 631 607 635
rect 611 631 612 635
rect 606 630 612 631
rect 608 613 610 630
rect 607 612 611 613
rect 607 607 611 608
rect 558 592 559 596
rect 563 592 564 596
rect 558 591 564 592
rect 570 595 576 596
rect 570 591 571 595
rect 575 591 576 595
rect 582 592 583 596
rect 587 592 588 596
rect 582 591 588 592
rect 594 595 600 596
rect 594 591 595 595
rect 599 591 600 595
rect 482 559 490 560
rect 482 555 483 559
rect 487 558 490 559
rect 550 563 556 564
rect 550 559 551 563
rect 555 559 556 563
rect 550 558 556 559
rect 487 555 488 558
rect 482 554 488 555
rect 484 532 486 554
rect 519 546 523 547
rect 519 541 523 542
rect 466 531 472 532
rect 466 527 467 531
rect 471 527 472 531
rect 466 526 472 527
rect 482 531 488 532
rect 482 527 483 531
rect 487 527 488 531
rect 482 526 488 527
rect 490 527 496 528
rect 468 488 470 526
rect 458 487 464 488
rect 458 483 459 487
rect 463 483 464 487
rect 458 482 464 483
rect 466 487 472 488
rect 466 483 467 487
rect 471 483 472 487
rect 466 482 472 483
rect 446 479 452 480
rect 446 475 447 479
rect 451 475 452 479
rect 446 474 452 475
rect 438 455 444 456
rect 438 451 439 455
rect 443 451 444 455
rect 438 450 444 451
rect 183 446 187 447
rect 183 441 187 442
rect 223 446 227 447
rect 230 446 236 447
rect 255 446 259 447
rect 223 441 227 442
rect 255 441 259 442
rect 279 446 283 447
rect 279 441 283 442
rect 303 446 307 447
rect 303 441 307 442
rect 327 446 331 447
rect 327 441 331 442
rect 343 446 347 447
rect 343 441 347 442
rect 379 446 383 447
rect 379 441 383 442
rect 447 446 451 447
rect 447 441 451 442
rect 184 417 186 441
rect 190 427 196 428
rect 190 423 191 427
rect 195 423 196 427
rect 190 422 196 423
rect 182 416 188 417
rect 182 412 183 416
rect 187 412 188 416
rect 182 411 188 412
rect 192 396 194 422
rect 224 419 226 441
rect 344 419 346 441
rect 222 418 228 419
rect 222 414 223 418
rect 227 414 228 418
rect 222 413 228 414
rect 342 418 348 419
rect 342 414 343 418
rect 347 414 348 418
rect 448 417 450 441
rect 342 413 348 414
rect 446 416 452 417
rect 446 412 447 416
rect 451 412 452 416
rect 446 411 452 412
rect 234 403 240 404
rect 234 399 235 403
rect 239 399 240 403
rect 234 398 240 399
rect 174 395 180 396
rect 174 391 175 395
rect 179 391 180 395
rect 174 390 180 391
rect 190 395 196 396
rect 190 391 191 395
rect 195 391 196 395
rect 190 390 196 391
rect 222 392 228 393
rect 192 387 194 390
rect 222 388 223 392
rect 227 388 228 392
rect 176 385 194 387
rect 206 387 212 388
rect 222 387 228 388
rect 158 384 164 385
rect 146 383 152 384
rect 134 382 140 383
rect 134 378 135 382
rect 139 378 140 382
rect 146 379 147 383
rect 151 379 152 383
rect 158 380 159 384
rect 163 380 164 384
rect 158 379 164 380
rect 146 378 152 379
rect 134 377 140 378
rect 136 355 138 377
rect 160 355 162 379
rect 111 354 115 355
rect 111 349 115 350
rect 135 354 139 355
rect 135 349 139 350
rect 159 354 163 355
rect 159 349 163 350
rect 112 298 114 349
rect 136 305 138 349
rect 150 327 156 328
rect 150 323 151 327
rect 155 323 156 327
rect 150 322 156 323
rect 134 304 140 305
rect 134 300 135 304
rect 139 300 140 304
rect 134 299 140 300
rect 110 297 116 298
rect 110 293 111 297
rect 115 293 116 297
rect 110 292 116 293
rect 110 279 116 280
rect 110 275 111 279
rect 115 275 116 279
rect 110 274 116 275
rect 112 243 114 274
rect 134 272 140 273
rect 134 268 135 272
rect 139 268 140 272
rect 134 267 140 268
rect 136 243 138 267
rect 111 242 115 243
rect 111 237 115 238
rect 135 242 139 243
rect 135 237 139 238
rect 143 242 147 243
rect 143 237 147 238
rect 112 218 114 237
rect 144 225 146 237
rect 142 224 148 225
rect 142 220 143 224
rect 147 220 148 224
rect 142 219 148 220
rect 110 217 116 218
rect 110 213 111 217
rect 115 213 116 217
rect 110 212 116 213
rect 152 204 154 322
rect 158 303 164 304
rect 158 299 159 303
rect 163 299 164 303
rect 158 298 164 299
rect 160 260 162 298
rect 176 260 178 385
rect 206 383 207 387
rect 211 386 212 387
rect 211 383 214 386
rect 182 382 188 383
rect 206 382 214 383
rect 182 378 183 382
rect 187 378 188 382
rect 182 377 188 378
rect 184 355 186 377
rect 212 372 214 382
rect 210 371 216 372
rect 210 367 211 371
rect 215 370 216 371
rect 215 367 218 370
rect 210 366 218 367
rect 194 359 200 360
rect 194 355 195 359
rect 199 355 200 359
rect 183 354 187 355
rect 194 354 200 355
rect 183 349 187 350
rect 184 297 186 349
rect 196 328 198 354
rect 206 351 212 352
rect 206 347 207 351
rect 211 347 212 351
rect 206 346 212 347
rect 208 328 210 346
rect 216 336 218 366
rect 224 355 226 387
rect 236 372 238 398
rect 342 392 348 393
rect 342 388 343 392
rect 347 388 348 392
rect 342 387 348 388
rect 426 387 432 388
rect 234 371 240 372
rect 234 367 235 371
rect 239 367 240 371
rect 234 366 240 367
rect 242 371 248 372
rect 242 367 243 371
rect 247 367 248 371
rect 242 366 248 367
rect 278 371 284 372
rect 278 367 279 371
rect 283 367 284 371
rect 278 366 284 367
rect 330 367 336 368
rect 223 354 227 355
rect 223 349 227 350
rect 214 335 220 336
rect 214 331 215 335
rect 219 331 220 335
rect 214 330 220 331
rect 194 327 200 328
rect 194 323 195 327
rect 199 323 200 327
rect 194 322 200 323
rect 206 327 212 328
rect 206 323 207 327
rect 211 323 212 327
rect 206 322 212 323
rect 182 296 188 297
rect 182 292 183 296
rect 187 292 188 296
rect 182 291 188 292
rect 208 288 210 322
rect 206 287 212 288
rect 206 283 207 287
rect 211 283 212 287
rect 206 282 212 283
rect 198 272 204 273
rect 198 268 199 272
rect 203 268 204 272
rect 198 267 204 268
rect 158 259 164 260
rect 158 255 159 259
rect 163 255 164 259
rect 158 254 164 255
rect 174 259 180 260
rect 174 255 175 259
rect 179 255 180 259
rect 174 254 180 255
rect 182 259 188 260
rect 182 255 183 259
rect 187 255 188 259
rect 182 254 188 255
rect 160 248 162 254
rect 158 247 164 248
rect 158 243 159 247
rect 163 243 164 247
rect 158 242 164 243
rect 167 242 171 243
rect 158 239 164 240
rect 158 235 159 239
rect 163 235 164 239
rect 167 237 171 238
rect 158 234 164 235
rect 150 203 156 204
rect 110 199 116 200
rect 110 195 111 199
rect 115 195 116 199
rect 150 199 151 203
rect 155 199 156 203
rect 150 198 156 199
rect 160 196 162 234
rect 168 225 170 237
rect 166 224 172 225
rect 166 220 167 224
rect 171 220 172 224
rect 166 219 172 220
rect 184 196 186 254
rect 200 243 202 267
rect 191 242 195 243
rect 191 237 195 238
rect 199 242 203 243
rect 199 237 203 238
rect 192 225 194 237
rect 208 232 210 282
rect 244 256 246 366
rect 280 364 302 366
rect 300 336 302 364
rect 330 363 331 367
rect 335 366 336 367
rect 335 363 338 366
rect 330 362 338 363
rect 322 359 328 360
rect 322 355 323 359
rect 327 355 328 359
rect 311 354 315 355
rect 322 354 328 355
rect 311 349 315 350
rect 286 335 292 336
rect 286 331 287 335
rect 291 331 292 335
rect 286 330 292 331
rect 298 335 304 336
rect 298 331 299 335
rect 303 331 304 335
rect 298 330 304 331
rect 270 327 276 328
rect 270 323 271 327
rect 275 323 276 327
rect 270 322 276 323
rect 242 255 248 256
rect 242 251 243 255
rect 247 251 248 255
rect 242 250 248 251
rect 244 240 246 250
rect 242 239 248 240
rect 242 235 243 239
rect 247 235 248 239
rect 242 234 248 235
rect 206 231 212 232
rect 206 227 207 231
rect 211 227 212 231
rect 206 226 212 227
rect 238 231 244 232
rect 238 227 239 231
rect 243 227 244 231
rect 238 226 244 227
rect 190 224 196 225
rect 190 220 191 224
rect 195 220 196 224
rect 190 219 196 220
rect 190 203 196 204
rect 190 199 191 203
rect 195 201 202 203
rect 195 199 196 201
rect 190 198 196 199
rect 110 194 116 195
rect 154 195 162 196
rect 112 135 114 194
rect 142 192 148 193
rect 142 188 143 192
rect 147 188 148 192
rect 154 191 155 195
rect 159 193 162 195
rect 178 195 186 196
rect 159 191 160 193
rect 154 190 160 191
rect 166 192 172 193
rect 142 187 148 188
rect 166 188 167 192
rect 171 188 172 192
rect 178 191 179 195
rect 183 193 186 195
rect 183 191 184 193
rect 178 190 184 191
rect 190 192 196 193
rect 166 187 172 188
rect 190 188 191 192
rect 195 188 196 192
rect 190 187 196 188
rect 200 192 202 201
rect 200 191 208 192
rect 200 187 203 191
rect 207 187 208 191
rect 144 135 146 187
rect 168 135 170 187
rect 192 135 194 187
rect 200 186 208 187
rect 210 187 216 188
rect 200 185 206 186
rect 204 164 206 185
rect 210 183 211 187
rect 215 183 216 187
rect 210 182 216 183
rect 218 187 224 188
rect 218 183 219 187
rect 223 183 224 187
rect 218 182 224 183
rect 202 163 208 164
rect 202 159 203 163
rect 207 159 208 163
rect 202 158 208 159
rect 212 140 214 182
rect 210 139 216 140
rect 210 135 211 139
rect 215 135 216 139
rect 111 134 115 135
rect 111 129 115 130
rect 135 134 139 135
rect 135 129 139 130
rect 143 134 147 135
rect 143 129 147 130
rect 167 134 171 135
rect 167 129 171 130
rect 191 134 195 135
rect 210 134 216 135
rect 191 129 195 130
rect 112 122 114 129
rect 134 128 140 129
rect 134 124 135 128
rect 139 124 140 128
rect 134 123 140 124
rect 110 121 116 122
rect 110 117 111 121
rect 115 117 116 121
rect 220 120 222 182
rect 240 148 242 226
rect 262 177 268 178
rect 262 173 263 177
rect 267 173 268 177
rect 262 172 268 173
rect 238 147 244 148
rect 238 143 239 147
rect 243 143 244 147
rect 238 142 244 143
rect 264 135 266 172
rect 272 164 274 322
rect 288 312 290 330
rect 286 311 292 312
rect 286 307 287 311
rect 291 307 292 311
rect 286 306 292 307
rect 312 297 314 349
rect 324 336 326 354
rect 322 335 328 336
rect 322 331 323 335
rect 327 334 328 335
rect 327 331 330 334
rect 322 330 330 331
rect 310 296 316 297
rect 310 292 311 296
rect 315 292 316 296
rect 310 291 316 292
rect 295 284 299 285
rect 295 279 299 280
rect 310 279 316 280
rect 296 260 298 279
rect 310 275 311 279
rect 315 275 316 279
rect 310 274 316 275
rect 294 259 300 260
rect 294 255 295 259
rect 299 255 300 259
rect 294 254 300 255
rect 302 251 308 252
rect 302 247 303 251
rect 307 247 308 251
rect 302 246 308 247
rect 279 242 283 243
rect 279 237 283 238
rect 280 224 282 237
rect 278 223 284 224
rect 278 219 279 223
rect 283 219 284 223
rect 278 218 284 219
rect 304 196 306 246
rect 312 243 314 274
rect 318 259 324 260
rect 318 255 319 259
rect 323 255 324 259
rect 318 254 324 255
rect 311 242 315 243
rect 311 237 315 238
rect 302 195 308 196
rect 302 191 303 195
rect 307 191 308 195
rect 302 190 308 191
rect 320 172 322 254
rect 318 171 324 172
rect 318 167 319 171
rect 323 167 324 171
rect 318 166 324 167
rect 328 164 330 330
rect 336 312 338 362
rect 344 355 346 387
rect 426 383 427 387
rect 431 383 432 387
rect 426 382 432 383
rect 446 384 452 385
rect 460 384 462 482
rect 484 467 486 526
rect 490 523 491 527
rect 495 523 496 527
rect 490 522 496 523
rect 492 480 494 522
rect 520 497 522 541
rect 552 520 554 558
rect 560 547 562 591
rect 570 590 576 591
rect 572 556 574 590
rect 570 555 576 556
rect 570 551 571 555
rect 575 551 576 555
rect 570 550 576 551
rect 584 547 586 591
rect 594 590 600 591
rect 559 546 563 547
rect 559 541 563 542
rect 575 546 579 547
rect 575 541 579 542
rect 583 546 587 547
rect 583 541 587 542
rect 550 519 556 520
rect 550 515 551 519
rect 555 515 556 519
rect 550 514 556 515
rect 518 496 524 497
rect 518 492 519 496
rect 523 492 524 496
rect 518 491 524 492
rect 576 489 578 541
rect 582 519 588 520
rect 582 515 583 519
rect 587 515 588 519
rect 582 514 588 515
rect 574 488 580 489
rect 574 484 575 488
rect 579 484 580 488
rect 574 483 580 484
rect 490 479 496 480
rect 490 475 491 479
rect 495 475 496 479
rect 490 474 496 475
rect 574 474 580 475
rect 574 470 575 474
rect 579 470 580 474
rect 574 469 580 470
rect 484 465 490 467
rect 471 446 475 447
rect 471 441 475 442
rect 472 417 474 441
rect 488 436 490 465
rect 518 464 524 465
rect 518 460 519 464
rect 523 460 524 464
rect 518 459 524 460
rect 520 447 522 459
rect 576 447 578 469
rect 584 456 586 514
rect 582 455 588 456
rect 582 451 583 455
rect 587 451 588 455
rect 582 450 588 451
rect 511 446 515 447
rect 511 441 515 442
rect 519 446 523 447
rect 519 441 523 442
rect 575 446 579 447
rect 575 441 579 442
rect 486 435 492 436
rect 486 431 487 435
rect 491 431 492 435
rect 486 430 492 431
rect 470 416 476 417
rect 470 412 471 416
rect 475 412 476 416
rect 470 411 476 412
rect 478 395 484 396
rect 478 391 479 395
rect 483 391 484 395
rect 478 390 484 391
rect 470 384 476 385
rect 343 354 347 355
rect 343 349 347 350
rect 415 354 419 355
rect 415 349 419 350
rect 334 311 340 312
rect 334 307 335 311
rect 339 307 340 311
rect 416 307 418 349
rect 334 306 340 307
rect 414 306 420 307
rect 336 172 338 306
rect 414 302 415 306
rect 419 302 420 306
rect 428 304 430 382
rect 446 380 447 384
rect 451 380 452 384
rect 446 379 452 380
rect 458 383 464 384
rect 458 379 459 383
rect 463 382 464 383
rect 463 379 466 382
rect 470 380 471 384
rect 475 380 476 384
rect 470 379 476 380
rect 448 355 450 379
rect 458 378 466 379
rect 454 371 460 372
rect 454 367 455 371
rect 459 367 460 371
rect 454 366 460 367
rect 439 354 443 355
rect 439 349 443 350
rect 447 354 451 355
rect 447 349 451 350
rect 440 305 442 349
rect 438 304 444 305
rect 414 301 420 302
rect 426 303 432 304
rect 426 298 427 303
rect 431 298 432 303
rect 438 300 439 304
rect 443 300 444 304
rect 438 299 444 300
rect 427 295 431 296
rect 422 291 428 292
rect 422 287 423 291
rect 427 287 428 291
rect 422 286 428 287
rect 414 272 420 273
rect 414 268 415 272
rect 419 268 420 272
rect 346 267 352 268
rect 414 267 420 268
rect 346 263 347 267
rect 351 263 352 267
rect 346 262 352 263
rect 334 171 340 172
rect 334 167 335 171
rect 339 167 340 171
rect 334 166 340 167
rect 270 163 276 164
rect 270 159 271 163
rect 275 159 276 163
rect 270 158 276 159
rect 326 163 332 164
rect 326 159 327 163
rect 331 159 332 163
rect 326 158 332 159
rect 272 148 274 158
rect 270 147 276 148
rect 270 143 271 147
rect 275 143 276 147
rect 270 142 276 143
rect 348 136 350 262
rect 416 243 418 267
rect 383 242 387 243
rect 383 237 387 238
rect 407 242 411 243
rect 407 237 411 238
rect 415 242 419 243
rect 415 237 419 238
rect 384 225 386 237
rect 390 235 396 236
rect 390 231 391 235
rect 395 231 396 235
rect 390 230 396 231
rect 382 224 388 225
rect 382 220 383 224
rect 387 220 388 224
rect 382 219 388 220
rect 392 212 394 230
rect 408 225 410 237
rect 406 224 412 225
rect 406 220 407 224
rect 411 220 412 224
rect 406 219 412 220
rect 390 211 396 212
rect 390 207 391 211
rect 395 207 396 211
rect 390 206 396 207
rect 382 192 388 193
rect 406 192 412 193
rect 382 188 383 192
rect 387 188 388 192
rect 382 187 388 188
rect 394 191 400 192
rect 394 187 395 191
rect 399 187 400 191
rect 406 188 407 192
rect 411 188 412 192
rect 406 187 412 188
rect 346 135 352 136
rect 384 135 386 187
rect 394 186 400 187
rect 396 148 398 186
rect 394 147 400 148
rect 394 143 395 147
rect 399 143 400 147
rect 394 142 400 143
rect 408 135 410 187
rect 424 144 426 286
rect 447 284 451 285
rect 446 279 447 284
rect 451 279 452 284
rect 446 278 452 279
rect 438 272 444 273
rect 438 268 439 272
rect 443 268 444 272
rect 438 267 444 268
rect 440 243 442 267
rect 456 248 458 366
rect 464 256 466 378
rect 472 355 474 379
rect 480 372 482 390
rect 488 372 490 430
rect 512 419 514 441
rect 554 427 560 428
rect 554 423 555 427
rect 559 423 560 427
rect 554 422 560 423
rect 510 418 516 419
rect 510 414 511 418
rect 515 414 516 418
rect 510 413 516 414
rect 510 392 516 393
rect 510 388 511 392
rect 515 388 516 392
rect 510 387 516 388
rect 478 371 484 372
rect 478 367 479 371
rect 483 367 484 371
rect 478 366 484 367
rect 486 371 492 372
rect 486 367 487 371
rect 491 367 492 371
rect 486 366 492 367
rect 512 355 514 387
rect 518 371 524 372
rect 518 367 519 371
rect 523 367 524 371
rect 518 366 524 367
rect 520 364 522 366
rect 518 363 524 364
rect 518 359 519 363
rect 523 359 524 363
rect 518 358 524 359
rect 471 354 475 355
rect 471 349 475 350
rect 503 354 507 355
rect 503 349 507 350
rect 511 354 515 355
rect 511 349 515 350
rect 490 327 496 328
rect 490 323 491 327
rect 495 323 496 327
rect 490 322 496 323
rect 492 313 494 322
rect 488 311 494 313
rect 488 272 490 311
rect 504 297 506 349
rect 520 348 522 358
rect 518 347 524 348
rect 518 343 519 347
rect 523 343 524 347
rect 518 342 524 343
rect 546 327 552 328
rect 546 323 547 327
rect 551 323 552 327
rect 546 322 552 323
rect 535 300 539 301
rect 502 296 508 297
rect 502 292 503 296
rect 507 292 508 296
rect 535 295 539 296
rect 494 291 500 292
rect 502 291 508 292
rect 494 287 495 291
rect 499 287 500 291
rect 494 286 500 287
rect 486 271 492 272
rect 486 267 487 271
rect 491 267 492 271
rect 486 266 492 267
rect 462 255 468 256
rect 462 251 463 255
rect 467 251 468 255
rect 462 250 468 251
rect 454 247 460 248
rect 454 243 455 247
rect 459 243 460 247
rect 486 247 492 248
rect 486 243 487 247
rect 491 243 492 247
rect 431 242 435 243
rect 431 237 435 238
rect 439 242 443 243
rect 454 242 460 243
rect 475 242 479 243
rect 486 242 492 243
rect 439 237 443 238
rect 475 237 479 238
rect 432 225 434 237
rect 466 235 472 236
rect 438 231 444 232
rect 438 227 439 231
rect 443 227 444 231
rect 466 231 467 235
rect 471 231 472 235
rect 466 230 472 231
rect 438 226 444 227
rect 430 224 436 225
rect 430 220 431 224
rect 435 220 436 224
rect 430 219 436 220
rect 430 192 436 193
rect 430 188 431 192
rect 435 188 436 192
rect 430 187 436 188
rect 422 143 428 144
rect 422 139 423 143
rect 427 139 428 143
rect 422 138 428 139
rect 432 135 434 187
rect 239 134 243 135
rect 239 129 243 130
rect 263 134 267 135
rect 346 131 347 135
rect 351 131 352 135
rect 346 130 352 131
rect 367 134 371 135
rect 263 129 267 130
rect 367 129 371 130
rect 383 134 387 135
rect 383 129 387 130
rect 407 134 411 135
rect 407 129 411 130
rect 431 134 435 135
rect 431 129 435 130
rect 238 128 244 129
rect 238 124 239 128
rect 243 124 244 128
rect 238 123 244 124
rect 366 128 372 129
rect 366 124 367 128
rect 371 124 372 128
rect 366 123 372 124
rect 110 116 116 117
rect 218 119 224 120
rect 218 115 219 119
rect 223 115 224 119
rect 440 116 442 226
rect 446 211 452 212
rect 446 207 447 211
rect 451 207 452 211
rect 446 206 452 207
rect 448 172 450 206
rect 468 204 470 230
rect 476 220 478 237
rect 474 219 480 220
rect 474 215 475 219
rect 479 215 480 219
rect 474 214 480 215
rect 454 203 460 204
rect 454 199 455 203
rect 459 199 460 203
rect 454 198 460 199
rect 466 203 472 204
rect 466 199 467 203
rect 471 199 472 203
rect 466 198 472 199
rect 474 200 480 201
rect 446 171 452 172
rect 446 167 447 171
rect 451 167 452 171
rect 446 166 452 167
rect 456 156 458 198
rect 474 196 475 200
rect 479 196 480 200
rect 474 195 480 196
rect 454 155 460 156
rect 454 151 455 155
rect 459 151 460 155
rect 454 150 460 151
rect 476 135 478 195
rect 488 156 490 242
rect 486 155 492 156
rect 486 151 487 155
rect 491 151 492 155
rect 486 150 492 151
rect 488 136 490 150
rect 496 148 498 286
rect 502 283 508 284
rect 502 279 503 283
rect 507 279 508 283
rect 502 278 508 279
rect 504 243 506 278
rect 503 242 507 243
rect 503 237 507 238
rect 536 208 538 295
rect 534 207 540 208
rect 534 203 535 207
rect 539 203 540 207
rect 534 202 540 203
rect 494 147 500 148
rect 494 143 495 147
rect 499 143 500 147
rect 494 142 500 143
rect 486 135 492 136
rect 475 134 479 135
rect 486 131 487 135
rect 491 131 492 135
rect 486 130 492 131
rect 495 134 499 135
rect 475 129 479 130
rect 495 129 499 130
rect 494 128 500 129
rect 494 124 495 128
rect 499 124 500 128
rect 494 123 500 124
rect 548 116 550 322
rect 556 264 558 422
rect 584 348 586 450
rect 596 372 598 590
rect 608 520 610 607
rect 620 579 622 638
rect 640 608 642 646
rect 648 618 650 653
rect 646 617 652 618
rect 646 613 647 617
rect 651 613 652 617
rect 646 612 652 613
rect 638 607 644 608
rect 638 603 639 607
rect 643 603 644 607
rect 638 602 644 603
rect 646 604 652 605
rect 646 600 647 604
rect 651 600 652 604
rect 646 599 652 600
rect 616 577 622 579
rect 616 540 618 577
rect 648 547 650 599
rect 672 576 674 662
rect 696 659 698 677
rect 695 658 699 659
rect 695 653 699 654
rect 678 643 684 644
rect 678 639 679 643
rect 683 639 684 643
rect 678 638 684 639
rect 670 575 676 576
rect 670 571 671 575
rect 675 571 676 575
rect 670 570 676 571
rect 647 546 651 547
rect 647 541 651 542
rect 614 539 620 540
rect 614 535 615 539
rect 619 535 620 539
rect 614 534 620 535
rect 606 519 612 520
rect 606 515 607 519
rect 611 515 612 519
rect 606 514 612 515
rect 608 428 610 514
rect 626 495 632 496
rect 626 491 627 495
rect 631 491 632 495
rect 626 490 632 491
rect 615 446 619 447
rect 615 441 619 442
rect 606 427 612 428
rect 606 423 607 427
rect 611 423 612 427
rect 606 422 612 423
rect 616 417 618 441
rect 614 416 620 417
rect 614 412 615 416
rect 619 412 620 416
rect 614 411 620 412
rect 606 395 612 396
rect 606 391 607 395
rect 611 391 612 395
rect 606 390 612 391
rect 594 371 600 372
rect 594 367 595 371
rect 599 367 600 371
rect 594 366 600 367
rect 582 347 588 348
rect 582 343 583 347
rect 587 343 588 347
rect 582 342 588 343
rect 554 263 560 264
rect 554 259 555 263
rect 559 259 560 263
rect 554 258 560 259
rect 566 255 572 256
rect 566 251 567 255
rect 571 251 572 255
rect 566 250 572 251
rect 568 236 570 250
rect 566 235 572 236
rect 566 231 567 235
rect 571 231 572 235
rect 566 230 572 231
rect 574 183 580 184
rect 574 179 575 183
rect 579 179 580 183
rect 574 178 580 179
rect 598 183 604 184
rect 598 179 599 183
rect 603 182 604 183
rect 608 182 610 390
rect 628 388 630 490
rect 680 488 682 638
rect 712 556 714 726
rect 710 555 716 556
rect 710 551 711 555
rect 715 551 716 555
rect 710 550 716 551
rect 703 546 707 547
rect 703 541 707 542
rect 686 503 692 504
rect 686 499 687 503
rect 691 499 692 503
rect 686 498 692 499
rect 678 487 684 488
rect 678 483 679 487
rect 683 483 684 487
rect 678 482 684 483
rect 655 446 659 447
rect 655 441 659 442
rect 656 419 658 441
rect 654 418 660 419
rect 654 414 655 418
rect 659 414 660 418
rect 654 413 660 414
rect 654 392 660 393
rect 654 388 655 392
rect 659 388 660 392
rect 626 387 632 388
rect 654 387 660 388
rect 614 384 620 385
rect 614 380 615 384
rect 619 380 620 384
rect 626 383 627 387
rect 631 383 632 387
rect 626 382 632 383
rect 614 379 620 380
rect 616 355 618 379
rect 646 359 652 360
rect 646 355 647 359
rect 651 355 652 359
rect 656 355 658 387
rect 688 372 690 498
rect 704 497 706 541
rect 712 504 714 550
rect 710 503 716 504
rect 710 499 711 503
rect 715 499 716 503
rect 710 498 716 499
rect 702 496 708 497
rect 702 492 703 496
rect 707 492 708 496
rect 702 491 708 492
rect 702 464 708 465
rect 702 460 703 464
rect 707 460 708 464
rect 702 459 708 460
rect 704 447 706 459
rect 703 446 707 447
rect 703 441 707 442
rect 714 439 720 440
rect 714 435 715 439
rect 719 435 720 439
rect 714 434 720 435
rect 698 431 704 432
rect 698 427 699 431
rect 703 427 704 431
rect 698 426 704 427
rect 686 371 692 372
rect 686 367 687 371
rect 691 367 692 371
rect 686 366 692 367
rect 666 355 672 356
rect 615 354 619 355
rect 615 349 619 350
rect 639 354 643 355
rect 646 354 652 355
rect 655 354 659 355
rect 639 349 643 350
rect 640 307 642 349
rect 648 347 650 354
rect 666 351 667 355
rect 671 351 672 355
rect 666 350 672 351
rect 679 354 683 355
rect 655 349 659 350
rect 648 345 654 347
rect 652 332 654 345
rect 658 339 664 340
rect 658 335 659 339
rect 663 335 664 339
rect 658 334 664 335
rect 650 331 656 332
rect 650 327 651 331
rect 655 327 656 331
rect 650 326 656 327
rect 652 308 654 326
rect 650 307 656 308
rect 638 306 644 307
rect 638 302 639 306
rect 643 302 644 306
rect 650 303 651 307
rect 655 303 656 307
rect 650 302 656 303
rect 638 301 644 302
rect 660 296 662 334
rect 668 324 670 350
rect 679 349 683 350
rect 666 323 672 324
rect 666 319 667 323
rect 671 319 672 323
rect 666 318 672 319
rect 680 297 682 349
rect 688 348 690 366
rect 686 347 692 348
rect 686 343 687 347
rect 691 343 692 347
rect 686 342 692 343
rect 688 324 690 342
rect 700 340 702 426
rect 716 368 718 434
rect 740 376 742 794
rect 760 676 762 962
rect 767 957 771 958
rect 823 962 827 963
rect 823 957 827 958
rect 768 921 770 957
rect 824 921 826 957
rect 766 920 772 921
rect 822 920 828 921
rect 836 920 838 990
rect 958 989 959 993
rect 963 989 964 993
rect 958 988 964 989
rect 938 987 944 988
rect 938 983 939 987
rect 943 983 944 987
rect 938 982 944 983
rect 940 972 942 982
rect 946 979 952 980
rect 946 975 947 979
rect 951 975 952 979
rect 946 974 952 975
rect 958 975 964 976
rect 938 971 944 972
rect 926 968 932 969
rect 926 964 927 968
rect 931 964 932 968
rect 938 967 939 971
rect 943 967 944 971
rect 938 966 944 967
rect 926 963 932 964
rect 887 962 891 963
rect 887 957 891 958
rect 927 962 931 963
rect 927 957 931 958
rect 888 921 890 957
rect 928 921 930 957
rect 886 920 892 921
rect 926 920 932 921
rect 948 920 950 974
rect 958 971 959 975
rect 963 971 964 975
rect 958 970 964 971
rect 960 963 962 970
rect 959 962 963 963
rect 959 957 963 958
rect 766 916 767 920
rect 771 916 772 920
rect 766 915 772 916
rect 814 919 820 920
rect 814 915 815 919
rect 819 915 820 919
rect 822 916 823 920
rect 827 916 828 920
rect 822 915 828 916
rect 834 919 840 920
rect 834 915 835 919
rect 839 915 840 919
rect 886 916 887 920
rect 891 916 892 920
rect 886 915 892 916
rect 918 919 924 920
rect 918 915 919 919
rect 923 915 924 919
rect 926 916 927 920
rect 931 916 932 920
rect 926 915 932 916
rect 946 919 952 920
rect 946 915 947 919
rect 951 915 952 919
rect 814 914 820 915
rect 834 914 840 915
rect 918 914 924 915
rect 946 914 952 915
rect 960 914 962 957
rect 766 888 772 889
rect 766 884 767 888
rect 771 884 772 888
rect 766 883 772 884
rect 768 871 770 883
rect 767 870 771 871
rect 767 865 771 866
rect 775 870 779 871
rect 775 865 779 866
rect 807 870 811 871
rect 807 865 811 866
rect 766 859 772 860
rect 766 855 767 859
rect 771 855 772 859
rect 766 854 772 855
rect 768 820 770 854
rect 776 841 778 865
rect 808 841 810 865
rect 816 859 818 914
rect 842 907 848 908
rect 842 903 843 907
rect 847 903 848 907
rect 842 902 848 903
rect 834 899 840 900
rect 834 895 835 899
rect 839 895 840 899
rect 834 894 840 895
rect 822 888 828 889
rect 822 884 823 888
rect 827 884 828 888
rect 822 883 828 884
rect 824 871 826 883
rect 823 870 827 871
rect 823 865 827 866
rect 816 857 830 859
rect 774 840 780 841
rect 774 836 775 840
rect 779 836 780 840
rect 774 835 780 836
rect 806 840 812 841
rect 806 836 807 840
rect 811 836 812 840
rect 806 835 812 836
rect 766 819 772 820
rect 766 815 767 819
rect 771 815 772 819
rect 766 814 772 815
rect 768 732 770 814
rect 828 812 830 857
rect 826 811 832 812
rect 774 808 780 809
rect 774 804 775 808
rect 779 804 780 808
rect 774 803 780 804
rect 806 808 812 809
rect 806 804 807 808
rect 811 804 812 808
rect 806 803 812 804
rect 818 807 824 808
rect 818 803 819 807
rect 823 803 824 807
rect 826 807 827 811
rect 831 807 832 811
rect 826 806 832 807
rect 776 759 778 803
rect 808 759 810 803
rect 818 802 824 803
rect 820 764 822 802
rect 836 796 838 894
rect 844 875 846 902
rect 886 888 892 889
rect 886 884 887 888
rect 891 884 892 888
rect 886 883 892 884
rect 840 873 846 875
rect 840 826 842 873
rect 888 871 890 883
rect 847 870 851 871
rect 847 865 851 866
rect 887 870 891 871
rect 887 865 891 866
rect 848 843 850 865
rect 898 851 904 852
rect 898 847 899 851
rect 903 847 904 851
rect 898 846 904 847
rect 846 842 852 843
rect 846 838 847 842
rect 851 838 852 842
rect 846 837 852 838
rect 840 824 858 826
rect 840 802 842 824
rect 846 816 852 817
rect 846 812 847 816
rect 851 812 852 816
rect 846 811 852 812
rect 840 800 846 802
rect 834 795 840 796
rect 834 791 835 795
rect 839 791 840 795
rect 834 790 840 791
rect 818 763 824 764
rect 836 763 838 790
rect 844 763 846 800
rect 818 759 819 763
rect 823 759 824 763
rect 775 758 779 759
rect 775 753 779 754
rect 799 758 803 759
rect 799 753 803 754
rect 807 758 811 759
rect 818 758 824 759
rect 828 761 838 763
rect 840 761 846 763
rect 828 755 830 761
rect 807 753 811 754
rect 824 753 830 755
rect 790 747 796 748
rect 790 743 791 747
rect 795 743 796 747
rect 790 742 796 743
rect 766 731 772 732
rect 766 727 767 731
rect 771 727 772 731
rect 766 726 772 727
rect 758 675 764 676
rect 758 671 759 675
rect 763 671 764 675
rect 758 670 764 671
rect 775 658 779 659
rect 775 653 779 654
rect 776 629 778 653
rect 774 628 780 629
rect 774 624 775 628
rect 779 624 780 628
rect 774 623 780 624
rect 782 607 788 608
rect 782 603 783 607
rect 787 603 788 607
rect 782 602 788 603
rect 774 596 780 597
rect 774 592 775 596
rect 779 592 780 596
rect 774 591 780 592
rect 776 547 778 591
rect 751 546 755 547
rect 751 541 755 542
rect 775 546 779 547
rect 775 541 779 542
rect 752 497 754 541
rect 784 528 786 602
rect 792 588 794 742
rect 800 717 802 753
rect 824 748 826 753
rect 840 752 842 761
rect 848 759 850 811
rect 856 796 858 824
rect 854 795 860 796
rect 854 791 855 795
rect 859 791 860 795
rect 854 790 860 791
rect 847 758 851 759
rect 847 753 851 754
rect 834 751 842 752
rect 822 747 828 748
rect 822 743 823 747
rect 827 743 828 747
rect 834 747 835 751
rect 839 748 842 751
rect 839 747 840 748
rect 834 746 840 747
rect 822 742 828 743
rect 798 716 804 717
rect 836 716 838 746
rect 798 712 799 716
rect 803 712 804 716
rect 798 711 804 712
rect 834 715 840 716
rect 834 711 835 715
rect 839 711 840 715
rect 834 710 840 711
rect 848 709 850 753
rect 858 747 864 748
rect 858 743 859 747
rect 863 743 864 747
rect 858 742 864 743
rect 866 747 872 748
rect 866 743 867 747
rect 871 743 872 747
rect 866 742 872 743
rect 846 708 852 709
rect 846 704 847 708
rect 851 704 852 708
rect 806 703 812 704
rect 846 703 852 704
rect 806 699 807 703
rect 811 699 812 703
rect 806 698 812 699
rect 798 684 804 685
rect 798 680 799 684
rect 803 680 804 684
rect 798 679 804 680
rect 800 659 802 679
rect 808 664 810 698
rect 846 691 852 692
rect 846 687 847 691
rect 851 687 852 691
rect 846 686 852 687
rect 834 671 840 672
rect 834 667 835 671
rect 839 667 840 671
rect 832 666 840 667
rect 832 665 838 666
rect 806 663 812 664
rect 806 659 807 663
rect 811 659 812 663
rect 799 658 803 659
rect 806 658 812 659
rect 818 663 824 664
rect 818 659 819 663
rect 823 659 824 663
rect 818 658 824 659
rect 799 653 803 654
rect 811 644 815 645
rect 810 639 811 644
rect 815 639 816 644
rect 810 638 816 639
rect 798 631 804 632
rect 798 627 799 631
rect 803 627 804 631
rect 798 626 804 627
rect 800 596 802 626
rect 798 595 804 596
rect 798 591 799 595
rect 803 591 804 595
rect 798 590 804 591
rect 790 587 796 588
rect 812 587 814 638
rect 820 611 822 658
rect 832 652 834 665
rect 848 659 850 686
rect 839 658 843 659
rect 839 653 843 654
rect 847 658 851 659
rect 847 653 851 654
rect 830 651 836 652
rect 830 647 831 651
rect 835 647 836 651
rect 830 646 836 647
rect 840 629 842 653
rect 838 628 844 629
rect 838 624 839 628
rect 843 624 844 628
rect 838 623 844 624
rect 790 583 791 587
rect 795 583 796 587
rect 790 582 796 583
rect 804 585 814 587
rect 816 609 822 611
rect 794 575 800 576
rect 794 571 795 575
rect 799 571 800 575
rect 794 570 800 571
rect 782 527 788 528
rect 762 523 768 524
rect 762 519 763 523
rect 767 519 768 523
rect 782 523 783 527
rect 787 523 788 527
rect 782 522 788 523
rect 762 518 768 519
rect 750 496 756 497
rect 764 496 766 518
rect 796 512 798 570
rect 794 511 800 512
rect 794 507 795 511
rect 799 507 800 511
rect 794 506 800 507
rect 750 492 751 496
rect 755 492 756 496
rect 750 491 756 492
rect 762 495 768 496
rect 762 491 763 495
rect 767 491 768 495
rect 804 494 806 585
rect 816 576 818 609
rect 822 604 828 605
rect 822 600 823 604
rect 827 600 828 604
rect 822 599 828 600
rect 814 575 820 576
rect 814 571 815 575
rect 819 571 820 575
rect 814 570 820 571
rect 810 563 816 564
rect 810 559 811 563
rect 815 559 816 563
rect 810 558 816 559
rect 812 508 814 558
rect 824 547 826 599
rect 846 575 852 576
rect 830 571 836 572
rect 830 567 831 571
rect 835 567 836 571
rect 846 571 847 575
rect 851 571 852 575
rect 846 570 852 571
rect 830 566 836 567
rect 832 556 834 566
rect 830 555 836 556
rect 830 551 831 555
rect 835 551 836 555
rect 830 550 836 551
rect 848 548 850 570
rect 846 547 852 548
rect 823 546 827 547
rect 823 541 827 542
rect 831 546 835 547
rect 846 543 847 547
rect 851 543 852 547
rect 846 542 852 543
rect 831 541 835 542
rect 832 512 834 541
rect 838 539 844 540
rect 838 535 839 539
rect 843 535 844 539
rect 838 534 844 535
rect 830 511 836 512
rect 810 507 816 508
rect 810 503 811 507
rect 815 503 816 507
rect 830 507 831 511
rect 835 507 836 511
rect 830 506 836 507
rect 810 502 816 503
rect 840 499 842 534
rect 762 490 768 491
rect 792 492 806 494
rect 828 497 842 499
rect 782 475 788 476
rect 782 471 783 475
rect 787 471 788 475
rect 782 470 788 471
rect 774 467 780 468
rect 750 464 756 465
rect 750 460 751 464
rect 755 460 756 464
rect 774 463 775 467
rect 779 463 780 467
rect 774 462 780 463
rect 763 460 767 461
rect 750 459 756 460
rect 752 447 754 459
rect 762 455 763 460
rect 767 455 768 460
rect 762 454 768 455
rect 766 447 772 448
rect 751 446 755 447
rect 766 443 767 447
rect 771 443 772 447
rect 766 442 772 443
rect 751 441 755 442
rect 738 375 744 376
rect 738 371 739 375
rect 743 371 744 375
rect 738 370 744 371
rect 714 367 720 368
rect 714 363 715 367
rect 719 363 720 367
rect 714 362 720 363
rect 698 339 704 340
rect 698 335 699 339
rect 703 335 704 339
rect 698 334 704 335
rect 700 324 702 334
rect 686 323 692 324
rect 686 319 687 323
rect 691 319 692 323
rect 686 318 692 319
rect 698 323 704 324
rect 698 319 699 323
rect 703 319 704 323
rect 698 318 704 319
rect 678 296 684 297
rect 658 295 664 296
rect 658 291 659 295
rect 663 291 664 295
rect 678 292 679 296
rect 683 292 684 296
rect 678 291 684 292
rect 658 290 664 291
rect 678 282 684 283
rect 678 278 679 282
rect 683 278 684 282
rect 678 277 684 278
rect 638 272 644 273
rect 638 268 639 272
rect 643 268 644 272
rect 638 267 644 268
rect 640 243 642 267
rect 646 263 652 264
rect 646 259 647 263
rect 651 259 652 263
rect 646 258 652 259
rect 623 242 627 243
rect 623 237 627 238
rect 639 242 643 243
rect 639 237 643 238
rect 624 215 626 237
rect 622 214 628 215
rect 622 210 623 214
rect 627 210 628 214
rect 622 209 628 210
rect 622 200 628 201
rect 622 196 623 200
rect 627 196 628 200
rect 622 195 628 196
rect 603 180 610 182
rect 603 179 604 180
rect 598 178 604 179
rect 576 156 578 178
rect 574 155 580 156
rect 574 151 575 155
rect 579 151 580 155
rect 574 150 580 151
rect 624 135 626 195
rect 634 191 640 192
rect 634 187 635 191
rect 639 187 640 191
rect 634 186 640 187
rect 623 134 627 135
rect 623 129 627 130
rect 622 128 628 129
rect 636 128 638 186
rect 648 172 650 258
rect 680 243 682 277
rect 679 242 683 243
rect 679 237 683 238
rect 642 171 650 172
rect 642 167 643 171
rect 647 168 650 171
rect 647 167 648 168
rect 642 166 648 167
rect 688 156 690 318
rect 716 184 718 362
rect 742 331 748 332
rect 742 327 743 331
rect 747 327 748 331
rect 742 326 748 327
rect 744 316 746 326
rect 742 315 748 316
rect 742 311 743 315
rect 747 311 748 315
rect 742 310 748 311
rect 768 308 770 442
rect 776 364 778 462
rect 784 440 786 470
rect 782 439 788 440
rect 782 435 783 439
rect 787 435 788 439
rect 782 434 788 435
rect 792 432 794 492
rect 799 446 803 447
rect 799 441 803 442
rect 790 431 796 432
rect 790 427 791 431
rect 795 427 796 431
rect 790 426 796 427
rect 792 424 794 426
rect 790 423 796 424
rect 790 419 791 423
rect 795 419 796 423
rect 790 418 796 419
rect 800 406 802 441
rect 828 440 830 497
rect 846 465 852 466
rect 846 461 847 465
rect 851 461 852 465
rect 846 460 852 461
rect 834 459 840 460
rect 834 455 835 459
rect 839 455 840 459
rect 834 454 840 455
rect 826 439 832 440
rect 826 435 827 439
rect 831 435 832 439
rect 826 434 832 435
rect 822 431 828 432
rect 822 427 823 431
rect 827 427 828 431
rect 822 426 828 427
rect 798 405 804 406
rect 798 401 799 405
rect 803 401 804 405
rect 798 400 804 401
rect 798 392 804 393
rect 798 388 799 392
rect 803 388 804 392
rect 798 387 804 388
rect 774 363 780 364
rect 774 359 775 363
rect 779 359 780 363
rect 774 358 780 359
rect 776 344 778 358
rect 800 355 802 387
rect 799 354 803 355
rect 799 349 803 350
rect 807 354 811 355
rect 807 349 811 350
rect 774 343 780 344
rect 774 339 775 343
rect 779 339 780 343
rect 774 338 780 339
rect 782 339 788 340
rect 766 307 772 308
rect 766 303 767 307
rect 771 303 772 307
rect 766 302 772 303
rect 776 260 778 338
rect 782 335 783 339
rect 787 335 788 339
rect 782 334 788 335
rect 774 259 780 260
rect 774 255 775 259
rect 779 255 780 259
rect 774 254 780 255
rect 742 247 748 248
rect 742 243 743 247
rect 747 243 748 247
rect 735 242 739 243
rect 742 242 748 243
rect 775 242 779 243
rect 735 237 739 238
rect 736 225 738 237
rect 734 224 740 225
rect 734 220 735 224
rect 739 220 740 224
rect 734 219 740 220
rect 744 204 746 242
rect 775 237 779 238
rect 776 225 778 237
rect 774 224 780 225
rect 774 220 775 224
rect 779 220 780 224
rect 774 219 780 220
rect 784 204 786 334
rect 808 296 810 349
rect 806 295 812 296
rect 806 291 807 295
rect 811 291 812 295
rect 806 290 812 291
rect 802 277 808 278
rect 802 273 803 277
rect 807 273 808 277
rect 802 272 808 273
rect 804 243 806 272
rect 803 242 807 243
rect 803 237 807 238
rect 815 242 819 243
rect 815 237 819 238
rect 816 225 818 237
rect 814 224 820 225
rect 814 220 815 224
rect 819 220 820 224
rect 814 219 820 220
rect 824 204 826 426
rect 836 364 838 454
rect 848 447 850 460
rect 860 448 862 742
rect 868 600 870 742
rect 900 645 902 846
rect 920 724 922 914
rect 958 913 964 914
rect 958 909 959 913
rect 963 909 964 913
rect 958 908 964 909
rect 946 907 952 908
rect 946 903 947 907
rect 951 903 952 907
rect 946 902 952 903
rect 926 888 932 889
rect 926 884 927 888
rect 931 884 932 888
rect 926 883 932 884
rect 928 871 930 883
rect 927 870 931 871
rect 927 865 931 866
rect 926 747 932 748
rect 926 743 927 747
rect 931 743 932 747
rect 926 742 932 743
rect 918 723 924 724
rect 918 719 919 723
rect 923 719 924 723
rect 918 718 924 719
rect 928 667 930 742
rect 938 679 944 680
rect 938 675 939 679
rect 943 675 944 679
rect 938 674 944 675
rect 920 665 930 667
rect 899 644 903 645
rect 899 639 903 640
rect 866 599 872 600
rect 866 595 867 599
rect 871 595 872 599
rect 866 594 872 595
rect 868 576 870 594
rect 866 575 872 576
rect 866 571 867 575
rect 871 571 872 575
rect 866 570 872 571
rect 878 571 884 572
rect 878 567 879 571
rect 883 567 884 571
rect 878 566 884 567
rect 870 555 876 556
rect 870 551 871 555
rect 875 551 876 555
rect 870 550 876 551
rect 872 524 874 550
rect 870 523 876 524
rect 870 519 871 523
rect 875 519 876 523
rect 870 518 876 519
rect 880 516 882 566
rect 906 531 912 532
rect 906 527 907 531
rect 911 527 912 531
rect 906 526 912 527
rect 908 523 910 526
rect 904 521 910 523
rect 878 515 884 516
rect 878 511 879 515
rect 883 514 884 515
rect 883 512 890 514
rect 883 511 884 512
rect 878 510 884 511
rect 870 499 876 500
rect 870 495 871 499
rect 875 495 876 499
rect 870 494 876 495
rect 872 448 874 494
rect 858 447 864 448
rect 847 446 851 447
rect 858 443 859 447
rect 863 443 864 447
rect 858 442 864 443
rect 870 447 876 448
rect 870 443 871 447
rect 875 443 876 447
rect 870 442 876 443
rect 847 441 851 442
rect 874 439 880 440
rect 874 435 875 439
rect 879 435 880 439
rect 874 434 880 435
rect 862 431 868 432
rect 862 427 863 431
rect 867 427 868 431
rect 862 426 868 427
rect 834 363 840 364
rect 834 359 835 363
rect 839 359 840 363
rect 834 358 840 359
rect 864 348 866 426
rect 862 347 868 348
rect 862 343 863 347
rect 867 343 868 347
rect 876 344 878 434
rect 862 342 868 343
rect 874 343 880 344
rect 830 339 836 340
rect 830 335 831 339
rect 835 335 836 339
rect 874 339 875 343
rect 879 339 880 343
rect 874 338 880 339
rect 830 334 836 335
rect 742 203 748 204
rect 742 199 743 203
rect 747 199 748 203
rect 742 198 748 199
rect 782 203 788 204
rect 782 199 783 203
rect 787 199 788 203
rect 782 198 788 199
rect 822 203 828 204
rect 822 199 823 203
rect 827 199 828 203
rect 822 198 828 199
rect 734 192 740 193
rect 774 192 780 193
rect 734 188 735 192
rect 739 188 740 192
rect 734 187 740 188
rect 746 191 752 192
rect 746 187 747 191
rect 751 187 752 191
rect 774 188 775 192
rect 779 188 780 192
rect 774 187 780 188
rect 814 192 820 193
rect 814 188 815 192
rect 819 188 820 192
rect 814 187 820 188
rect 714 183 720 184
rect 714 179 715 183
rect 719 179 720 183
rect 714 178 720 179
rect 686 155 692 156
rect 686 151 687 155
rect 691 151 692 155
rect 686 150 692 151
rect 736 135 738 187
rect 746 186 752 187
rect 748 176 750 186
rect 758 183 764 184
rect 758 179 759 183
rect 763 179 764 183
rect 758 178 764 179
rect 746 175 752 176
rect 746 171 747 175
rect 751 171 752 175
rect 746 170 752 171
rect 748 156 750 170
rect 746 155 752 156
rect 746 151 747 155
rect 751 151 752 155
rect 746 150 752 151
rect 735 134 739 135
rect 735 129 739 130
rect 751 134 755 135
rect 751 129 755 130
rect 750 128 756 129
rect 622 124 623 128
rect 627 124 628 128
rect 622 123 628 124
rect 634 127 640 128
rect 634 123 635 127
rect 639 123 640 127
rect 750 124 751 128
rect 755 124 756 128
rect 750 123 756 124
rect 634 122 640 123
rect 760 116 762 178
rect 776 135 778 187
rect 816 135 818 187
rect 832 184 834 334
rect 862 323 868 324
rect 862 319 863 323
rect 867 319 868 323
rect 862 318 868 319
rect 864 292 866 318
rect 878 307 884 308
rect 878 303 879 307
rect 883 303 884 307
rect 878 302 884 303
rect 862 291 868 292
rect 862 287 863 291
rect 867 287 868 291
rect 862 286 868 287
rect 855 242 859 243
rect 855 237 859 238
rect 856 225 858 237
rect 854 224 860 225
rect 854 220 855 224
rect 859 220 860 224
rect 854 219 860 220
rect 854 192 860 193
rect 880 192 882 302
rect 888 204 890 512
rect 904 340 906 521
rect 920 507 922 665
rect 927 658 931 659
rect 927 653 931 654
rect 928 629 930 653
rect 926 628 932 629
rect 926 624 927 628
rect 931 624 932 628
rect 926 623 932 624
rect 926 596 932 597
rect 940 596 942 674
rect 926 592 927 596
rect 931 592 932 596
rect 926 591 932 592
rect 938 595 944 596
rect 938 591 939 595
rect 943 591 944 595
rect 928 547 930 591
rect 938 590 944 591
rect 927 546 931 547
rect 927 541 931 542
rect 940 531 942 590
rect 948 564 950 902
rect 958 895 964 896
rect 958 891 959 895
rect 963 891 964 895
rect 958 890 964 891
rect 960 871 962 890
rect 959 870 963 871
rect 959 865 963 866
rect 960 834 962 865
rect 958 833 964 834
rect 958 829 959 833
rect 963 829 964 833
rect 958 828 964 829
rect 958 815 964 816
rect 958 811 959 815
rect 963 811 964 815
rect 958 810 964 811
rect 960 759 962 810
rect 959 758 963 759
rect 959 753 963 754
rect 960 710 962 753
rect 958 709 964 710
rect 958 705 959 709
rect 963 705 964 709
rect 958 704 964 705
rect 958 691 964 692
rect 958 687 959 691
rect 963 687 964 691
rect 958 686 964 687
rect 960 659 962 686
rect 959 658 963 659
rect 959 653 963 654
rect 960 622 962 653
rect 958 621 964 622
rect 958 617 959 621
rect 963 617 964 621
rect 958 616 964 617
rect 958 603 964 604
rect 958 599 959 603
rect 963 599 964 603
rect 958 598 964 599
rect 946 563 952 564
rect 946 559 947 563
rect 951 559 952 563
rect 946 558 952 559
rect 960 547 962 598
rect 959 546 963 547
rect 959 541 963 542
rect 916 505 922 507
rect 936 529 942 531
rect 916 482 918 505
rect 912 480 918 482
rect 910 479 916 480
rect 910 475 911 479
rect 915 475 916 479
rect 910 474 916 475
rect 910 455 916 456
rect 910 451 911 455
rect 915 451 916 455
rect 910 450 916 451
rect 912 356 914 450
rect 918 447 924 448
rect 918 443 919 447
rect 923 443 924 447
rect 918 442 924 443
rect 927 446 931 447
rect 920 404 922 442
rect 927 441 931 442
rect 928 417 930 441
rect 926 416 932 417
rect 926 412 927 416
rect 931 412 932 416
rect 926 411 932 412
rect 918 403 924 404
rect 918 399 919 403
rect 923 399 924 403
rect 918 398 924 399
rect 910 355 916 356
rect 910 351 911 355
rect 915 351 916 355
rect 910 350 916 351
rect 902 339 908 340
rect 902 335 903 339
rect 907 335 908 339
rect 902 334 908 335
rect 904 316 906 334
rect 902 315 908 316
rect 902 311 903 315
rect 907 311 908 315
rect 902 310 908 311
rect 903 242 907 243
rect 903 237 907 238
rect 904 225 906 237
rect 902 224 908 225
rect 902 220 903 224
rect 907 220 908 224
rect 902 219 908 220
rect 912 204 914 350
rect 920 312 922 398
rect 936 396 938 529
rect 960 490 962 541
rect 958 489 964 490
rect 958 485 959 489
rect 963 485 964 489
rect 958 484 964 485
rect 958 471 964 472
rect 958 467 959 471
rect 963 467 964 471
rect 958 466 964 467
rect 960 447 962 466
rect 959 446 963 447
rect 959 441 963 442
rect 960 410 962 441
rect 958 409 964 410
rect 958 405 959 409
rect 963 405 964 409
rect 958 404 964 405
rect 934 395 940 396
rect 934 391 935 395
rect 939 391 940 395
rect 934 390 940 391
rect 958 391 964 392
rect 926 384 932 385
rect 926 380 927 384
rect 931 380 932 384
rect 926 379 932 380
rect 928 355 930 379
rect 927 354 931 355
rect 927 349 931 350
rect 918 311 924 312
rect 918 307 919 311
rect 923 307 924 311
rect 918 306 924 307
rect 928 305 930 349
rect 936 348 938 390
rect 958 387 959 391
rect 963 387 964 391
rect 958 386 964 387
rect 960 355 962 386
rect 959 354 963 355
rect 959 349 963 350
rect 934 347 940 348
rect 934 343 935 347
rect 939 343 940 347
rect 934 342 940 343
rect 926 304 932 305
rect 926 300 927 304
rect 931 300 932 304
rect 926 299 932 300
rect 960 298 962 349
rect 958 297 964 298
rect 958 293 959 297
rect 963 293 964 297
rect 958 292 964 293
rect 946 291 952 292
rect 946 287 947 291
rect 951 287 952 291
rect 946 286 952 287
rect 926 272 932 273
rect 926 268 927 272
rect 931 268 932 272
rect 926 267 932 268
rect 928 243 930 267
rect 934 259 940 260
rect 934 255 935 259
rect 939 255 940 259
rect 934 254 940 255
rect 927 242 931 243
rect 927 237 931 238
rect 928 225 930 237
rect 926 224 932 225
rect 926 220 927 224
rect 931 220 932 224
rect 926 219 932 220
rect 936 204 938 254
rect 886 203 892 204
rect 886 199 887 203
rect 891 199 892 203
rect 886 198 892 199
rect 910 203 916 204
rect 910 199 911 203
rect 915 199 916 203
rect 910 198 916 199
rect 934 203 940 204
rect 934 199 935 203
rect 939 199 940 203
rect 934 198 940 199
rect 854 188 855 192
rect 859 188 860 192
rect 854 187 860 188
rect 878 191 884 192
rect 878 187 879 191
rect 883 187 884 191
rect 830 183 836 184
rect 830 179 831 183
rect 835 179 836 183
rect 830 178 836 179
rect 856 135 858 187
rect 878 186 884 187
rect 888 184 890 198
rect 902 192 908 193
rect 948 192 950 286
rect 958 279 964 280
rect 958 275 959 279
rect 963 275 964 279
rect 958 274 964 275
rect 960 243 962 274
rect 959 242 963 243
rect 959 237 963 238
rect 960 218 962 237
rect 958 217 964 218
rect 958 213 959 217
rect 963 213 964 217
rect 958 212 964 213
rect 958 199 964 200
rect 958 195 959 199
rect 963 195 964 199
rect 958 194 964 195
rect 902 188 903 192
rect 907 188 908 192
rect 946 191 952 192
rect 902 187 908 188
rect 926 190 932 191
rect 886 183 892 184
rect 886 179 887 183
rect 891 179 892 183
rect 886 178 892 179
rect 904 135 906 187
rect 926 186 927 190
rect 931 186 932 190
rect 946 187 947 191
rect 951 187 952 191
rect 946 186 952 187
rect 926 185 932 186
rect 928 135 930 185
rect 960 135 962 194
rect 775 134 779 135
rect 775 129 779 130
rect 815 134 819 135
rect 815 129 819 130
rect 855 134 859 135
rect 855 129 859 130
rect 903 134 907 135
rect 903 129 907 130
rect 927 134 931 135
rect 927 129 931 130
rect 959 134 963 135
rect 959 129 963 130
rect 960 122 962 129
rect 958 121 964 122
rect 958 117 959 121
rect 963 117 964 121
rect 958 116 964 117
rect 218 114 224 115
rect 438 115 444 116
rect 438 111 439 115
rect 443 111 444 115
rect 438 110 444 111
rect 546 115 552 116
rect 546 111 547 115
rect 551 111 552 115
rect 546 110 552 111
rect 758 115 764 116
rect 758 111 759 115
rect 763 111 764 115
rect 758 110 764 111
rect 110 103 116 104
rect 110 99 111 103
rect 115 99 116 103
rect 110 98 116 99
rect 958 103 964 104
rect 958 99 959 103
rect 963 99 964 103
rect 958 98 964 99
rect 112 91 114 98
rect 134 96 140 97
rect 134 92 135 96
rect 139 92 140 96
rect 134 91 140 92
rect 238 96 244 97
rect 238 92 239 96
rect 243 92 244 96
rect 238 91 244 92
rect 366 96 372 97
rect 366 92 367 96
rect 371 92 372 96
rect 366 91 372 92
rect 494 96 500 97
rect 494 92 495 96
rect 499 92 500 96
rect 494 91 500 92
rect 622 96 628 97
rect 622 92 623 96
rect 627 92 628 96
rect 622 91 628 92
rect 750 96 756 97
rect 750 92 751 96
rect 755 92 756 96
rect 750 91 756 92
rect 960 91 962 98
rect 111 90 115 91
rect 111 85 115 86
rect 135 90 139 91
rect 135 85 139 86
rect 239 90 243 91
rect 239 85 243 86
rect 367 90 371 91
rect 367 85 371 86
rect 495 90 499 91
rect 495 85 499 86
rect 623 90 627 91
rect 623 85 627 86
rect 751 90 755 91
rect 751 85 755 86
rect 959 90 963 91
rect 959 85 963 86
<< m4c >>
rect 111 1002 115 1006
rect 135 1002 139 1006
rect 319 1002 323 1006
rect 527 1002 531 1006
rect 735 1002 739 1006
rect 927 1002 931 1006
rect 959 1002 963 1006
rect 111 958 115 962
rect 135 958 139 962
rect 159 958 163 962
rect 183 958 187 962
rect 111 866 115 870
rect 135 866 139 870
rect 159 866 163 870
rect 111 754 115 758
rect 135 754 139 758
rect 175 866 179 870
rect 183 866 187 870
rect 231 958 235 962
rect 311 958 315 962
rect 319 958 323 962
rect 231 866 235 870
rect 159 754 163 758
rect 175 754 179 758
rect 455 958 459 962
rect 519 958 523 962
rect 527 958 531 962
rect 583 958 587 962
rect 647 958 651 962
rect 711 958 715 962
rect 735 958 739 962
rect 311 866 315 870
rect 279 754 283 758
rect 111 654 115 658
rect 135 654 139 658
rect 159 654 163 658
rect 175 654 179 658
rect 111 542 115 546
rect 327 866 331 870
rect 303 754 307 758
rect 311 754 315 758
rect 327 754 331 758
rect 351 754 355 758
rect 451 866 455 870
rect 459 866 463 870
rect 383 754 387 758
rect 415 754 419 758
rect 439 754 443 758
rect 451 754 455 758
rect 463 754 467 758
rect 279 654 283 658
rect 151 542 155 546
rect 159 542 163 546
rect 111 442 115 446
rect 135 442 139 446
rect 151 442 155 446
rect 159 442 163 446
rect 275 611 279 612
rect 275 608 279 611
rect 303 654 307 658
rect 327 654 331 658
rect 351 654 355 658
rect 383 654 387 658
rect 255 542 259 546
rect 279 542 283 546
rect 287 542 291 546
rect 303 542 307 546
rect 327 542 331 546
rect 379 542 383 546
rect 415 654 419 658
rect 439 654 443 658
rect 439 542 443 546
rect 455 654 459 658
rect 463 654 467 658
rect 519 866 523 870
rect 575 866 579 870
rect 583 866 587 870
rect 495 754 499 758
rect 543 754 547 758
rect 587 792 591 796
rect 575 754 579 758
rect 639 866 643 870
rect 647 866 651 870
rect 639 754 643 758
rect 655 754 659 758
rect 711 866 715 870
rect 695 754 699 758
rect 495 654 499 658
rect 543 654 547 658
rect 559 654 563 658
rect 583 654 587 658
rect 647 654 651 658
rect 655 654 659 658
rect 607 608 611 612
rect 519 542 523 546
rect 183 442 187 446
rect 223 442 227 446
rect 255 442 259 446
rect 279 442 283 446
rect 303 442 307 446
rect 327 442 331 446
rect 343 442 347 446
rect 379 442 383 446
rect 447 442 451 446
rect 111 350 115 354
rect 135 350 139 354
rect 159 350 163 354
rect 111 238 115 242
rect 135 238 139 242
rect 143 238 147 242
rect 183 350 187 354
rect 223 350 227 354
rect 167 238 171 242
rect 191 238 195 242
rect 199 238 203 242
rect 311 350 315 354
rect 111 130 115 134
rect 135 130 139 134
rect 143 130 147 134
rect 167 130 171 134
rect 191 130 195 134
rect 295 280 299 284
rect 279 238 283 242
rect 311 238 315 242
rect 559 542 563 546
rect 575 542 579 546
rect 583 542 587 546
rect 471 442 475 446
rect 511 442 515 446
rect 519 442 523 446
rect 575 442 579 446
rect 343 350 347 354
rect 415 350 419 354
rect 439 350 443 354
rect 447 350 451 354
rect 427 299 431 300
rect 427 296 431 299
rect 383 238 387 242
rect 407 238 411 242
rect 415 238 419 242
rect 447 283 451 284
rect 447 280 451 283
rect 471 350 475 354
rect 503 350 507 354
rect 511 350 515 354
rect 535 296 539 300
rect 431 238 435 242
rect 439 238 443 242
rect 475 238 479 242
rect 239 130 243 134
rect 263 130 267 134
rect 367 130 371 134
rect 383 130 387 134
rect 407 130 411 134
rect 431 130 435 134
rect 503 238 507 242
rect 475 130 479 134
rect 495 130 499 134
rect 695 654 699 658
rect 647 542 651 546
rect 615 442 619 446
rect 703 542 707 546
rect 655 442 659 446
rect 703 442 707 446
rect 615 350 619 354
rect 639 350 643 354
rect 655 350 659 354
rect 679 350 683 354
rect 767 958 771 962
rect 823 958 827 962
rect 887 958 891 962
rect 927 958 931 962
rect 959 958 963 962
rect 767 866 771 870
rect 775 866 779 870
rect 807 866 811 870
rect 823 866 827 870
rect 847 866 851 870
rect 887 866 891 870
rect 775 754 779 758
rect 799 754 803 758
rect 807 754 811 758
rect 775 654 779 658
rect 751 542 755 546
rect 775 542 779 546
rect 847 754 851 758
rect 799 654 803 658
rect 811 643 815 644
rect 811 640 815 643
rect 839 654 843 658
rect 847 654 851 658
rect 823 542 827 546
rect 831 542 835 546
rect 763 459 767 460
rect 763 456 767 459
rect 751 442 755 446
rect 623 238 627 242
rect 639 238 643 242
rect 623 130 627 134
rect 679 238 683 242
rect 799 442 803 446
rect 799 350 803 354
rect 807 350 811 354
rect 735 238 739 242
rect 775 238 779 242
rect 803 238 807 242
rect 815 238 819 242
rect 927 866 931 870
rect 899 640 903 644
rect 847 442 851 446
rect 735 130 739 134
rect 751 130 755 134
rect 855 238 859 242
rect 927 654 931 658
rect 927 542 931 546
rect 959 866 963 870
rect 959 754 963 758
rect 959 654 963 658
rect 959 542 963 546
rect 927 442 931 446
rect 903 238 907 242
rect 959 442 963 446
rect 927 350 931 354
rect 959 350 963 354
rect 927 238 931 242
rect 959 238 963 242
rect 775 130 779 134
rect 815 130 819 134
rect 855 130 859 134
rect 903 130 907 134
rect 927 130 931 134
rect 959 130 963 134
rect 111 86 115 90
rect 135 86 139 90
rect 239 86 243 90
rect 367 86 371 90
rect 495 86 499 90
rect 623 86 627 90
rect 751 86 755 90
rect 959 86 963 90
<< m4 >>
rect 84 1001 85 1007
rect 91 1006 983 1007
rect 91 1002 111 1006
rect 115 1002 135 1006
rect 139 1002 319 1006
rect 323 1002 527 1006
rect 531 1002 735 1006
rect 739 1002 927 1006
rect 931 1002 959 1006
rect 963 1002 983 1006
rect 91 1001 983 1002
rect 989 1001 990 1007
rect 96 957 97 963
rect 103 962 995 963
rect 103 958 111 962
rect 115 958 135 962
rect 139 958 159 962
rect 163 958 183 962
rect 187 958 231 962
rect 235 958 311 962
rect 315 958 319 962
rect 323 958 455 962
rect 459 958 519 962
rect 523 958 527 962
rect 531 958 583 962
rect 587 958 647 962
rect 651 958 711 962
rect 715 958 735 962
rect 739 958 767 962
rect 771 958 823 962
rect 827 958 887 962
rect 891 958 927 962
rect 931 958 959 962
rect 963 958 995 962
rect 103 957 995 958
rect 1001 957 1002 963
rect 84 865 85 871
rect 91 870 983 871
rect 91 866 111 870
rect 115 866 135 870
rect 139 866 159 870
rect 163 866 175 870
rect 179 866 183 870
rect 187 866 231 870
rect 235 866 311 870
rect 315 866 327 870
rect 331 866 451 870
rect 455 866 459 870
rect 463 866 519 870
rect 523 866 575 870
rect 579 866 583 870
rect 587 866 639 870
rect 643 866 647 870
rect 651 866 711 870
rect 715 866 767 870
rect 771 866 775 870
rect 779 866 807 870
rect 811 866 823 870
rect 827 866 847 870
rect 851 866 887 870
rect 891 866 927 870
rect 931 866 959 870
rect 963 866 983 870
rect 91 865 983 866
rect 989 865 990 871
rect 586 796 592 797
rect 638 796 639 797
rect 586 792 587 796
rect 591 792 639 796
rect 586 791 592 792
rect 638 791 639 792
rect 645 791 646 797
rect 96 753 97 759
rect 103 758 995 759
rect 103 754 111 758
rect 115 754 135 758
rect 139 754 159 758
rect 163 754 175 758
rect 179 754 279 758
rect 283 754 303 758
rect 307 754 311 758
rect 315 754 327 758
rect 331 754 351 758
rect 355 754 383 758
rect 387 754 415 758
rect 419 754 439 758
rect 443 754 451 758
rect 455 754 463 758
rect 467 754 495 758
rect 499 754 543 758
rect 547 754 575 758
rect 579 754 639 758
rect 643 754 655 758
rect 659 754 695 758
rect 699 754 775 758
rect 779 754 799 758
rect 803 754 807 758
rect 811 754 847 758
rect 851 754 959 758
rect 963 754 995 758
rect 103 753 995 754
rect 1001 753 1002 759
rect 84 653 85 659
rect 91 658 983 659
rect 91 654 111 658
rect 115 654 135 658
rect 139 654 159 658
rect 163 654 175 658
rect 179 654 279 658
rect 283 654 303 658
rect 307 654 327 658
rect 331 654 351 658
rect 355 654 383 658
rect 387 654 415 658
rect 419 654 439 658
rect 443 654 455 658
rect 459 654 463 658
rect 467 654 495 658
rect 499 654 543 658
rect 547 654 559 658
rect 563 654 583 658
rect 587 654 647 658
rect 651 654 655 658
rect 659 654 695 658
rect 699 654 775 658
rect 779 654 799 658
rect 803 654 839 658
rect 843 654 847 658
rect 851 654 927 658
rect 931 654 959 658
rect 963 654 983 658
rect 91 653 983 654
rect 989 653 990 659
rect 810 644 816 645
rect 898 644 904 645
rect 810 640 811 644
rect 815 640 899 644
rect 903 640 904 644
rect 810 639 816 640
rect 898 639 904 640
rect 274 612 280 613
rect 606 612 612 613
rect 274 608 275 612
rect 279 608 607 612
rect 611 608 612 612
rect 274 607 280 608
rect 606 607 612 608
rect 96 541 97 547
rect 103 546 995 547
rect 103 542 111 546
rect 115 542 151 546
rect 155 542 159 546
rect 163 542 255 546
rect 259 542 279 546
rect 283 542 287 546
rect 291 542 303 546
rect 307 542 327 546
rect 331 542 379 546
rect 383 542 439 546
rect 443 542 519 546
rect 523 542 559 546
rect 563 542 575 546
rect 579 542 583 546
rect 587 542 647 546
rect 651 542 703 546
rect 707 542 751 546
rect 755 542 775 546
rect 779 542 823 546
rect 827 542 831 546
rect 835 542 927 546
rect 931 542 959 546
rect 963 542 995 546
rect 103 541 995 542
rect 1001 541 1002 547
rect 638 455 639 461
rect 645 460 646 461
rect 762 460 768 461
rect 645 456 763 460
rect 767 456 768 460
rect 645 455 646 456
rect 762 455 768 456
rect 84 441 85 447
rect 91 446 983 447
rect 91 442 111 446
rect 115 442 135 446
rect 139 442 151 446
rect 155 442 159 446
rect 163 442 183 446
rect 187 442 223 446
rect 227 442 255 446
rect 259 442 279 446
rect 283 442 303 446
rect 307 442 327 446
rect 331 442 343 446
rect 347 442 379 446
rect 383 442 447 446
rect 451 442 471 446
rect 475 442 511 446
rect 515 442 519 446
rect 523 442 575 446
rect 579 442 615 446
rect 619 442 655 446
rect 659 442 703 446
rect 707 442 751 446
rect 755 442 799 446
rect 803 442 847 446
rect 851 442 927 446
rect 931 442 959 446
rect 963 442 983 446
rect 91 441 983 442
rect 989 441 990 447
rect 96 349 97 355
rect 103 354 995 355
rect 103 350 111 354
rect 115 350 135 354
rect 139 350 159 354
rect 163 350 183 354
rect 187 350 223 354
rect 227 350 311 354
rect 315 350 343 354
rect 347 350 415 354
rect 419 350 439 354
rect 443 350 447 354
rect 451 350 471 354
rect 475 350 503 354
rect 507 350 511 354
rect 515 350 615 354
rect 619 350 639 354
rect 643 350 655 354
rect 659 350 679 354
rect 683 350 799 354
rect 803 350 807 354
rect 811 350 927 354
rect 931 350 959 354
rect 963 350 995 354
rect 103 349 995 350
rect 1001 349 1002 355
rect 426 300 432 301
rect 534 300 540 301
rect 426 296 427 300
rect 431 296 535 300
rect 539 296 540 300
rect 426 295 432 296
rect 534 295 540 296
rect 294 284 300 285
rect 446 284 452 285
rect 294 280 295 284
rect 299 280 447 284
rect 451 280 452 284
rect 294 279 300 280
rect 446 279 452 280
rect 84 237 85 243
rect 91 242 983 243
rect 91 238 111 242
rect 115 238 135 242
rect 139 238 143 242
rect 147 238 167 242
rect 171 238 191 242
rect 195 238 199 242
rect 203 238 279 242
rect 283 238 311 242
rect 315 238 383 242
rect 387 238 407 242
rect 411 238 415 242
rect 419 238 431 242
rect 435 238 439 242
rect 443 238 475 242
rect 479 238 503 242
rect 507 238 623 242
rect 627 238 639 242
rect 643 238 679 242
rect 683 238 735 242
rect 739 238 775 242
rect 779 238 803 242
rect 807 238 815 242
rect 819 238 855 242
rect 859 238 903 242
rect 907 238 927 242
rect 931 238 959 242
rect 963 238 983 242
rect 91 237 983 238
rect 989 237 990 243
rect 96 129 97 135
rect 103 134 995 135
rect 103 130 111 134
rect 115 130 135 134
rect 139 130 143 134
rect 147 130 167 134
rect 171 130 191 134
rect 195 130 239 134
rect 243 130 263 134
rect 267 130 367 134
rect 371 130 383 134
rect 387 130 407 134
rect 411 130 431 134
rect 435 130 475 134
rect 479 130 495 134
rect 499 130 623 134
rect 627 130 735 134
rect 739 130 751 134
rect 755 130 775 134
rect 779 130 815 134
rect 819 130 855 134
rect 859 130 903 134
rect 907 130 927 134
rect 931 130 959 134
rect 963 130 995 134
rect 103 129 995 130
rect 1001 129 1002 135
rect 84 85 85 91
rect 91 90 983 91
rect 91 86 111 90
rect 115 86 135 90
rect 139 86 239 90
rect 243 86 367 90
rect 371 86 495 90
rect 499 86 623 90
rect 627 86 751 90
rect 755 86 959 90
rect 963 86 983 90
rect 91 85 983 86
rect 989 85 990 91
<< m5c >>
rect 85 1001 91 1007
rect 983 1001 989 1007
rect 97 957 103 963
rect 995 957 1001 963
rect 85 865 91 871
rect 983 865 989 871
rect 639 791 645 797
rect 97 753 103 759
rect 995 753 1001 759
rect 85 653 91 659
rect 983 653 989 659
rect 97 541 103 547
rect 995 541 1001 547
rect 639 455 645 461
rect 85 441 91 447
rect 983 441 989 447
rect 97 349 103 355
rect 995 349 1001 355
rect 85 237 91 243
rect 983 237 989 243
rect 97 129 103 135
rect 995 129 1001 135
rect 85 85 91 91
rect 983 85 989 91
<< m5 >>
rect 84 1007 92 1008
rect 84 1001 85 1007
rect 91 1001 92 1007
rect 84 871 92 1001
rect 84 865 85 871
rect 91 865 92 871
rect 84 659 92 865
rect 84 653 85 659
rect 91 653 92 659
rect 84 447 92 653
rect 84 441 85 447
rect 91 441 92 447
rect 84 243 92 441
rect 84 237 85 243
rect 91 237 92 243
rect 84 91 92 237
rect 84 85 85 91
rect 91 85 92 91
rect 84 72 92 85
rect 96 963 104 1008
rect 96 957 97 963
rect 103 957 104 963
rect 96 759 104 957
rect 982 1007 990 1008
rect 982 1001 983 1007
rect 989 1001 990 1007
rect 982 871 990 1001
rect 982 865 983 871
rect 989 865 990 871
rect 638 797 646 798
rect 638 791 639 797
rect 645 791 646 797
rect 638 790 646 791
rect 96 753 97 759
rect 103 753 104 759
rect 96 547 104 753
rect 96 541 97 547
rect 103 541 104 547
rect 96 355 104 541
rect 640 462 644 790
rect 982 659 990 865
rect 982 653 983 659
rect 989 653 990 659
rect 638 461 646 462
rect 638 455 639 461
rect 645 455 646 461
rect 638 454 646 455
rect 96 349 97 355
rect 103 349 104 355
rect 96 135 104 349
rect 96 129 97 135
rect 103 129 104 135
rect 96 72 104 129
rect 982 447 990 653
rect 982 441 983 447
rect 989 441 990 447
rect 982 243 990 441
rect 982 237 983 243
rect 989 237 990 243
rect 982 91 990 237
rect 982 85 983 91
rect 989 85 990 91
rect 982 72 990 85
rect 994 963 1002 1008
rect 994 957 995 963
rect 1001 957 1002 963
rect 994 759 1002 957
rect 994 753 995 759
rect 1001 753 1002 759
rect 994 547 1002 753
rect 994 541 995 547
rect 1001 541 1002 547
rect 994 355 1002 541
rect 994 349 995 355
rect 1001 349 1002 355
rect 994 135 1002 349
rect 994 129 995 135
rect 1001 129 1002 135
rect 994 72 1002 129
use welltap_svt  __well_tap__0
timestamp 1753821931
transform 1 0 104 0 1 96
box 8 4 12 24
use welltap_svt  __well_tap__1
timestamp 1753821931
transform 1 0 952 0 1 96
box 8 4 12 24
use welltap_svt  __well_tap__2
timestamp 1753821931
transform 1 0 104 0 -1 220
box 8 4 12 24
use welltap_svt  __well_tap__3
timestamp 1753821931
transform 1 0 952 0 -1 220
box 8 4 12 24
use welltap_svt  __well_tap__4
timestamp 1753821931
transform 1 0 104 0 1 272
box 8 4 12 24
use welltap_svt  __well_tap__5
timestamp 1753821931
transform 1 0 952 0 1 272
box 8 4 12 24
use welltap_svt  __well_tap__6
timestamp 1753821931
transform 1 0 104 0 -1 412
box 8 4 12 24
use welltap_svt  __well_tap__7
timestamp 1753821931
transform 1 0 952 0 -1 412
box 8 4 12 24
use welltap_svt  __well_tap__8
timestamp 1753821931
transform 1 0 104 0 1 464
box 8 4 12 24
use welltap_svt  __well_tap__9
timestamp 1753821931
transform 1 0 952 0 1 464
box 8 4 12 24
use welltap_svt  __well_tap__10
timestamp 1753821931
transform 1 0 104 0 -1 624
box 8 4 12 24
use welltap_svt  __well_tap__11
timestamp 1753821931
transform 1 0 952 0 -1 624
box 8 4 12 24
use welltap_svt  __well_tap__12
timestamp 1753821931
transform 1 0 104 0 1 684
box 8 4 12 24
use welltap_svt  __well_tap__13
timestamp 1753821931
transform 1 0 952 0 1 684
box 8 4 12 24
use welltap_svt  __well_tap__14
timestamp 1753821931
transform 1 0 104 0 -1 836
box 8 4 12 24
use welltap_svt  __well_tap__15
timestamp 1753821931
transform 1 0 952 0 -1 836
box 8 4 12 24
use welltap_svt  __well_tap__16
timestamp 1753821931
transform 1 0 104 0 1 888
box 8 4 12 24
use welltap_svt  __well_tap__17
timestamp 1753821931
transform 1 0 952 0 1 888
box 8 4 12 24
use welltap_svt  __well_tap__18
timestamp 1753821931
transform 1 0 104 0 -1 996
box 8 4 12 24
use welltap_svt  __well_tap__19
timestamp 1753821931
transform 1 0 952 0 -1 996
box 8 4 12 24
use _0_0cell_0_0ginvx0  c_aB_acx0 ~/Desktop/Testing_for_Learning/Layout/post_layout/mag2ext/test
timestamp 1753821931
transform 1 0 488 0 1 88
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aB_acx1
timestamp 1753821931
transform 1 0 616 0 1 88
box 5 4 23 41
use _0_0cell_0_0g0n1n2n3naaa_02ox0  c_aC_50_6_acx0 ~/Desktop/Testing_for_Learning/Layout/post_layout/mag2ext/test
timestamp 1753821931
transform 1 0 656 0 1 260
box 5 4 116 67
use _0_0cell_0_0g0n1n2n3naaa_04256aaaox0  c_aC_50_6_acx1 ~/Desktop/Testing_for_Learning/Layout/post_layout/mag2ext/test
timestamp 1753821931
transform 1 0 792 0 -1 648
box 8 3 123 80
use _0_0cell_0_0g0n1n2na3n2n4n5naaa2n6n7naaooa_082a92aoox0  c_aC_50_6_acx2 ~/Desktop/Testing_for_Learning/Layout/post_layout/mag2ext/test
timestamp 1753821931
transform 1 0 776 0 1 444
box 5 5 161 98
use _0_0cell_0_0g0n1n2n3n4naaaa_0536aaox0  c_aC_50_6_acx3 ~/Desktop/Testing_for_Learning/Layout/post_layout/mag2ext/test
timestamp 1753821931
transform 1 0 816 0 1 664
box 5 2 123 87
use _0_0cell_0_0g0n1n2n3n4n5naaaaa_0653aaox0  c_aC_50_6_acx4 ~/Desktop/Testing_for_Learning/Layout/post_layout/mag2ext/test
timestamp 1753821931
transform 1 0 776 0 1 260
box 5 3 139 88
use _0_0cell_0_0g0n1n2n3n4naaao_025a4267aaooax0  c_aC_50_6_acx5 ~/Desktop/Testing_for_Learning/Layout/post_layout/mag2ext/test
timestamp 1753821931
transform 1 0 752 0 -1 444
box 8 4 161 88
use _0_0cell_0_0g0n1n2naa_032aox0  c_aC_50_6_acx6 ~/Desktop/Testing_for_Learning/Layout/post_layout/mag2ext/test
timestamp 1753821931
transform 1 0 824 0 -1 856
box 5 5 117 68
use _0_0cell_0_0g0n1n2naa_032aox0  c_aC_50_6_acx7
timestamp 1753821931
transform 1 0 632 0 -1 432
box 5 5 117 68
use _0_0cell_0_0ginvx0  c_aC_50_6_acx8
timestamp 1753821931
transform 1 0 920 0 1 880
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_50_6_acx9
timestamp 1753821931
transform 1 0 808 0 -1 228
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_50_6_acx10
timestamp 1753821931
transform 1 0 768 0 -1 632
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_50_6_acx11
timestamp 1753821931
transform 1 0 744 0 1 456
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_50_6_acx12
timestamp 1753821931
transform 1 0 848 0 -1 228
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_50_6_acx13
timestamp 1753821931
transform 1 0 896 0 -1 228
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_50_6_acx14
timestamp 1753821931
transform 1 0 920 0 -1 420
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_50_6_acx15
timestamp 1753821931
transform 1 0 920 0 -1 632
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_50_6_acx16
timestamp 1753821931
transform 1 0 816 0 1 880
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_50_6_acx17
timestamp 1753821931
transform 1 0 792 0 1 676
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_50_6_acx18
timestamp 1753821931
transform 1 0 744 0 1 88
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_50_6_acx19
timestamp 1753821931
transform 1 0 768 0 -1 228
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_50_6_acx20
timestamp 1753821931
transform 1 0 880 0 1 880
box 5 4 23 41
use _0_0cell_0_0ginvx1  c_aC_50_6_acx21 ~/Desktop/Testing_for_Learning/Layout/post_layout/mag2ext/test
timestamp 1753821931
transform 1 0 632 0 1 264
box 5 4 23 43
use _0_0cell_0_0ginvx0  c_aC_50_6_acx22
timestamp 1753821931
transform 1 0 920 0 1 264
box 5 4 23 41
use _0_0cell_0_0ginvx1  c_aC_50_6_acx23
timestamp 1753821931
transform 1 0 920 0 -1 228
box 5 4 23 43
use _0_0cell_0_0g0n1n2n3naaa_02ox0  c_aC_51_6_acx0
timestamp 1753821931
transform 1 0 520 0 1 672
box 5 4 116 67
use _0_0cell_0_0g0n1n2n3naaa_04256aaaox0  c_aC_51_6_acx1
timestamp 1753821931
transform 1 0 128 0 -1 860
box 8 3 123 80
use _0_0cell_0_0g0n1n2na3n2n4n5naaa2n6n7naaooa_082a92aoox0  c_aC_51_6_acx2
timestamp 1753821931
transform 1 0 256 0 -1 856
box 5 5 161 98
use _0_0cell_0_0g0n1n2n3n4naaaa_0536aaox0  c_aC_51_6_acx3
timestamp 1753821931
transform 1 0 280 0 1 868
box 5 2 123 87
use _0_0cell_0_0g0n1n2n3n4n5naaaaa_0653aaox0  c_aC_51_6_acx4
timestamp 1753821931
transform 1 0 424 0 -1 848
box 5 3 139 88
use _0_0cell_0_0g0n1n2n3n4naaao_025a4267aaooax0  c_aC_51_6_acx5
timestamp 1753821931
transform 1 0 592 0 -1 868
box 8 4 161 88
use _0_0cell_0_0g0n1n2naa_032aox0  c_aC_51_6_acx6
timestamp 1753821931
transform 1 0 152 0 1 664
box 5 5 117 68
use _0_0cell_0_0g0n1n2naa_032aox0  c_aC_51_6_acx7
timestamp 1753821931
transform 1 0 672 0 1 664
box 5 5 117 68
use _0_0cell_0_0ginvx0  c_aC_51_6_acx8
timestamp 1753821931
transform 1 0 128 0 -1 1004
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_51_6_acx9
timestamp 1753821931
transform 1 0 640 0 1 880
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_51_6_acx10
timestamp 1753821931
transform 1 0 152 0 1 880
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_51_6_acx11
timestamp 1753821931
transform 1 0 224 0 1 880
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_51_6_acx12
timestamp 1753821931
transform 1 0 448 0 1 880
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_51_6_acx13
timestamp 1753821931
transform 1 0 512 0 1 880
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_51_6_acx14
timestamp 1753821931
transform 1 0 576 0 1 880
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_51_6_acx15
timestamp 1753821931
transform 1 0 128 0 1 880
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_51_6_acx16
timestamp 1753821931
transform 1 0 760 0 1 880
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_51_6_acx17
timestamp 1753821931
transform 1 0 176 0 1 880
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_51_6_acx18
timestamp 1753821931
transform 1 0 768 0 -1 844
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_51_6_acx19
timestamp 1753821931
transform 1 0 704 0 1 880
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_51_6_acx20
timestamp 1753821931
transform 1 0 800 0 -1 844
box 5 4 23 41
use _0_0cell_0_0ginvx1  c_aC_51_6_acx21
timestamp 1753821931
transform 1 0 344 0 1 676
box 5 4 23 43
use _0_0cell_0_0ginvx0  c_aC_51_6_acx22
timestamp 1753821931
transform 1 0 568 0 -1 844
box 5 4 23 41
use _0_0cell_0_0ginvx1  c_aC_51_6_acx23
timestamp 1753821931
transform 1 0 488 0 1 676
box 5 4 23 43
use _0_0cell_0_0g0n1n2n3naaa_02ox0  c_aC_52_6_acx0
timestamp 1753821931
transform 1 0 552 0 1 452
box 5 4 116 67
use _0_0cell_0_0g0n1n2n3naaa_04256aaaox0  c_aC_52_6_acx1
timestamp 1753821931
transform 1 0 256 0 -1 648
box 8 3 123 80
use _0_0cell_0_0g0n1n2na3n2n4n5naaa2n6n7naaooa_082a92aoox0  c_aC_52_6_acx2
timestamp 1753821931
transform 1 0 384 0 -1 644
box 5 5 161 98
use _0_0cell_0_0g0n1n2n3n4naaaa_0536aaox0  c_aC_52_6_acx3
timestamp 1753821931
transform 1 0 128 0 -1 644
box 5 2 123 87
use _0_0cell_0_0g0n1n2n3n4n5naaaaa_0653aaox0  c_aC_52_6_acx4
timestamp 1753821931
transform 1 0 352 0 1 452
box 5 3 139 88
use _0_0cell_0_0g0n1n2n3n4naaao_025a4267aaooax0  c_aC_52_6_acx5
timestamp 1753821931
transform 1 0 600 0 -1 656
box 8 4 161 88
use _0_0cell_0_0g0n1n2naa_032aox0  c_aC_52_6_acx6
timestamp 1753821931
transform 1 0 128 0 1 444
box 5 5 117 68
use _0_0cell_0_0g0n1n2naa_032aox0  c_aC_52_6_acx7
timestamp 1753821931
transform 1 0 488 0 -1 432
box 5 5 117 68
use _0_0cell_0_0ginvx0  c_aC_52_6_acx8
timestamp 1753821931
transform 1 0 296 0 1 456
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_52_6_acx9
timestamp 1753821931
transform 1 0 696 0 1 456
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_52_6_acx10
timestamp 1753821931
transform 1 0 320 0 1 676
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_52_6_acx11
timestamp 1753821931
transform 1 0 376 0 1 676
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_52_6_acx12
timestamp 1753821931
transform 1 0 320 0 1 456
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_52_6_acx13
timestamp 1753821931
transform 1 0 552 0 -1 632
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_52_6_acx14
timestamp 1753821931
transform 1 0 512 0 1 456
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_52_6_acx15
timestamp 1753821931
transform 1 0 272 0 1 676
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_52_6_acx16
timestamp 1753821931
transform 1 0 128 0 1 676
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_52_6_acx17
timestamp 1753821931
transform 1 0 296 0 1 676
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_52_6_acx18
timestamp 1753821931
transform 1 0 648 0 1 676
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_52_6_acx19
timestamp 1753821931
transform 1 0 576 0 -1 632
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_52_6_acx20
timestamp 1753821931
transform 1 0 456 0 1 676
box 5 4 23 41
use _0_0cell_0_0ginvx1  c_aC_52_6_acx21
timestamp 1753821931
transform 1 0 128 0 -1 420
box 5 4 23 43
use _0_0cell_0_0ginvx0  c_aC_52_6_acx22
timestamp 1753821931
transform 1 0 432 0 1 676
box 5 4 23 41
use _0_0cell_0_0ginvx1  c_aC_52_6_acx23
timestamp 1753821931
transform 1 0 408 0 1 676
box 5 4 23 43
use _0_0cell_0_0g0n1n2n3naaa_02ox0  c_aC_53_6_acx0
timestamp 1753821931
transform 1 0 600 0 -1 232
box 5 4 116 67
use _0_0cell_0_0g0n1n2n3naaa_04256aaaox0  c_aC_53_6_acx1
timestamp 1753821931
transform 1 0 152 0 1 248
box 8 3 123 80
use _0_0cell_0_0g0n1n2na3n2n4n5naaa2n6n7naaooa_082a92aoox0  c_aC_53_6_acx2
timestamp 1753821931
transform 1 0 208 0 -1 240
box 5 5 161 98
use _0_0cell_0_0g0n1n2n3n4naaaa_0536aaox0  c_aC_53_6_acx3
timestamp 1753821931
transform 1 0 280 0 1 252
box 5 2 123 87
use _0_0cell_0_0g0n1n2n3n4n5naaaaa_0653aaox0  c_aC_53_6_acx4
timestamp 1753821931
transform 1 0 448 0 -1 232
box 5 3 139 88
use _0_0cell_0_0g0n1n2n3n4naaao_025a4267aaooax0  c_aC_53_6_acx5
timestamp 1753821931
transform 1 0 456 0 1 240
box 8 4 161 88
use _0_0cell_0_0g0n1n2naa_032aox0  c_aC_53_6_acx6
timestamp 1753821931
transform 1 0 200 0 -1 432
box 5 5 117 68
use _0_0cell_0_0g0n1n2naa_032aox0  c_aC_53_6_acx7
timestamp 1753821931
transform 1 0 320 0 -1 432
box 5 5 117 68
use _0_0cell_0_0ginvx0  c_aC_53_6_acx8
timestamp 1753821931
transform 1 0 128 0 1 88
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_53_6_acx9
timestamp 1753821931
transform 1 0 728 0 -1 228
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_53_6_acx10
timestamp 1753821931
transform 1 0 160 0 -1 228
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_53_6_acx11
timestamp 1753821931
transform 1 0 184 0 -1 228
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_53_6_acx12
timestamp 1753821931
transform 1 0 400 0 -1 228
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_53_6_acx13
timestamp 1753821931
transform 1 0 376 0 -1 228
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_53_6_acx14
timestamp 1753821931
transform 1 0 432 0 1 264
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_53_6_acx15
timestamp 1753821931
transform 1 0 128 0 1 264
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_53_6_acx16
timestamp 1753821931
transform 1 0 152 0 -1 420
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_53_6_acx17
timestamp 1753821931
transform 1 0 136 0 -1 228
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_53_6_acx18
timestamp 1753821931
transform 1 0 464 0 -1 420
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_53_6_acx19
timestamp 1753821931
transform 1 0 424 0 -1 228
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aC_53_6_acx20
timestamp 1753821931
transform 1 0 608 0 -1 420
box 5 4 23 41
use _0_0cell_0_0ginvx1  c_aC_53_6_acx21
timestamp 1753821931
transform 1 0 176 0 -1 420
box 5 4 23 43
use _0_0cell_0_0ginvx0  c_aC_53_6_acx22
timestamp 1753821931
transform 1 0 440 0 -1 420
box 5 4 23 41
use _0_0cell_0_0ginvx1  c_aC_53_6_acx23
timestamp 1753821931
transform 1 0 408 0 1 264
box 5 4 23 43
use _0_0cell_0_0ginvx0  c_aR_50_6_acx0
timestamp 1753821931
transform 1 0 920 0 -1 1004
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aR_50_6_acx1
timestamp 1753821931
transform 1 0 728 0 -1 1004
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aR_51_6_acx0
timestamp 1753821931
transform 1 0 312 0 -1 1004
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aR_51_6_acx1
timestamp 1753821931
transform 1 0 520 0 -1 1004
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aR_52_6_acx0
timestamp 1753821931
transform 1 0 272 0 1 456
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aR_52_6_acx1
timestamp 1753821931
transform 1 0 248 0 1 456
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aR_53_6_acx0
timestamp 1753821931
transform 1 0 232 0 1 88
box 5 4 23 41
use _0_0cell_0_0ginvx0  c_aR_53_6_acx1
timestamp 1753821931
transform 1 0 360 0 1 88
box 5 4 23 41
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
<< labels >>
flabel m1 s 550 1004 554 1008 0 FreeSans 24 0 0 0 IN.d[0]
port 0 nsew signal input
flabel m1 s 550 72 554 76 0 FreeSans 24 0 0 0 IN.d[1]
port 1 nsew signal input
flabel m1 s 1012 694 1016 698 0 FreeSans 24 0 0 0 IN.r
port 2 nsew signal input
flabel m1 s 1012 382 1016 386 0 FreeSans 24 0 0 0 IN.a
port 3 nsew signal output
flabel m1 s 80 538 84 542 0 FreeSans 24 0 0 0 Reset
port 4 nsew signal input
<< properties >>
string FIXED_BBOX 80 72 1016 1008
<< end >>
