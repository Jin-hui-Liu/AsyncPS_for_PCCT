magic
tech sky130A
magscale 1 2
timestamp 1753381912
<< nwell >>
rect 75 615 510 1140
rect 75 555 660 615
rect 75 375 1185 555
rect 1440 375 2085 1140
<< nmos >>
rect 375 210 405 300
rect 480 210 540 300
rect 780 210 810 300
rect 855 210 1185 300
rect 1290 75 1320 300
rect 1665 75 1695 300
rect 1935 75 1965 300
<< pmos >>
rect 195 420 225 1095
rect 270 420 300 1095
rect 375 420 405 1095
rect 480 420 540 570
rect 780 420 810 510
rect 855 420 1065 510
rect 1560 420 1590 1095
rect 1665 420 1695 1095
rect 1935 420 1965 1095
<< ndiff >>
rect 300 285 375 300
rect 300 240 315 285
rect 360 240 375 285
rect 300 210 375 240
rect 405 285 480 300
rect 405 240 420 285
rect 465 240 480 285
rect 405 210 480 240
rect 540 285 615 300
rect 540 240 555 285
rect 600 240 615 285
rect 540 210 615 240
rect 705 285 780 300
rect 705 240 720 285
rect 765 240 780 285
rect 705 210 780 240
rect 810 210 855 300
rect 1185 285 1290 300
rect 1185 240 1215 285
rect 1260 240 1290 285
rect 1185 210 1290 240
rect 1230 75 1290 210
rect 1320 150 1395 300
rect 1320 105 1335 150
rect 1380 105 1395 150
rect 1320 75 1395 105
rect 1590 285 1665 300
rect 1590 240 1605 285
rect 1650 240 1665 285
rect 1590 75 1665 240
rect 1695 270 1770 300
rect 1695 225 1710 270
rect 1755 225 1770 270
rect 1695 75 1770 225
rect 1860 270 1935 300
rect 1860 225 1875 270
rect 1920 225 1935 270
rect 1860 75 1935 225
rect 1965 150 2040 300
rect 1965 105 1980 150
rect 2025 105 2040 150
rect 1965 75 2040 105
<< pdiff >>
rect 120 1065 195 1095
rect 120 1020 135 1065
rect 180 1020 195 1065
rect 120 420 195 1020
rect 225 420 270 1095
rect 300 420 375 1095
rect 405 570 465 1095
rect 1485 990 1560 1095
rect 1485 945 1500 990
rect 1545 945 1560 990
rect 405 495 480 570
rect 405 450 420 495
rect 465 450 480 495
rect 405 420 480 450
rect 540 480 615 570
rect 540 435 555 480
rect 600 435 615 480
rect 540 420 615 435
rect 705 480 780 510
rect 705 435 720 480
rect 765 435 780 480
rect 705 420 780 435
rect 810 420 855 510
rect 1065 495 1140 510
rect 1065 450 1080 495
rect 1125 450 1140 495
rect 1065 420 1140 450
rect 1485 420 1560 945
rect 1590 420 1665 1095
rect 1695 1065 1770 1095
rect 1695 1020 1710 1065
rect 1755 1020 1770 1065
rect 1695 420 1770 1020
rect 1860 675 1935 1095
rect 1860 630 1875 675
rect 1920 630 1935 675
rect 1860 420 1935 630
rect 1965 990 2040 1095
rect 1965 945 1980 990
rect 2025 945 2040 990
rect 1965 420 2040 945
<< ndiffc >>
rect 315 240 360 285
rect 420 240 465 285
rect 555 240 600 285
rect 720 240 765 285
rect 1215 240 1260 285
rect 1335 105 1380 150
rect 1605 240 1650 285
rect 1710 225 1755 270
rect 1875 225 1920 270
rect 1980 105 2025 150
<< pdiffc >>
rect 135 1020 180 1065
rect 1500 945 1545 990
rect 420 450 465 495
rect 555 435 600 480
rect 720 435 765 480
rect 1080 450 1125 495
rect 1710 1020 1755 1065
rect 1875 630 1920 675
rect 1980 945 2025 990
<< poly >>
rect 240 1290 345 1320
rect 240 1245 270 1290
rect 315 1245 345 1290
rect 90 1215 195 1245
rect 240 1215 345 1245
rect 90 1170 120 1215
rect 165 1170 195 1215
rect 90 1140 225 1170
rect 195 1095 225 1140
rect 270 1095 300 1215
rect 405 1200 510 1230
rect 405 1155 435 1200
rect 480 1155 510 1200
rect 375 1125 510 1155
rect 1485 1215 1590 1245
rect 1485 1170 1515 1215
rect 1560 1170 1590 1215
rect 1485 1140 1590 1170
rect 375 1095 405 1125
rect 1560 1095 1590 1140
rect 1665 1215 1770 1245
rect 1665 1170 1695 1215
rect 1740 1170 1770 1215
rect 1665 1140 1770 1170
rect 1905 1200 2010 1230
rect 1905 1155 1935 1200
rect 1980 1155 2010 1200
rect 1665 1095 1695 1140
rect 1905 1125 2010 1155
rect 1935 1095 1965 1125
rect 480 675 615 705
rect 480 630 540 675
rect 585 630 615 675
rect 480 600 615 630
rect 930 615 1035 645
rect 480 570 540 600
rect 930 570 960 615
rect 1005 570 1035 615
rect 930 540 1035 570
rect 780 510 810 540
rect 855 510 1065 540
rect 1290 420 1395 450
rect 195 390 225 420
rect 270 390 300 420
rect 375 300 405 420
rect 480 300 540 420
rect 780 300 810 420
rect 855 390 1065 420
rect 1290 375 1320 420
rect 1365 375 1395 420
rect 1560 390 1590 420
rect 1290 345 1395 375
rect 855 300 1185 330
rect 1290 300 1320 345
rect 1665 300 1695 420
rect 1935 300 1965 420
rect 375 180 405 210
rect 480 180 540 210
rect 780 165 810 210
rect 855 180 1185 210
rect 705 135 810 165
rect 705 90 735 135
rect 780 90 810 135
rect 705 60 810 90
rect 1065 150 1170 180
rect 1065 105 1095 150
rect 1140 105 1170 150
rect 1065 75 1170 105
rect 1290 45 1320 75
rect 1665 45 1695 75
rect 1935 45 1965 75
<< polycont >>
rect 270 1245 315 1290
rect 120 1170 165 1215
rect 435 1155 480 1200
rect 1515 1170 1560 1215
rect 1695 1170 1740 1215
rect 1935 1155 1980 1200
rect 540 630 585 675
rect 960 570 1005 615
rect 1320 375 1365 420
rect 735 90 780 135
rect 1095 105 1140 150
<< locali >>
rect 240 1290 345 1320
rect 240 1245 270 1290
rect 315 1245 345 1290
rect 90 1215 195 1245
rect 240 1215 345 1245
rect 90 1170 120 1215
rect 165 1170 195 1215
rect 90 1140 195 1170
rect 405 1200 510 1230
rect 405 1155 435 1200
rect 480 1155 510 1200
rect 405 1125 510 1155
rect 1485 1215 1590 1245
rect 1485 1170 1515 1215
rect 1560 1170 1590 1215
rect 1485 1140 1590 1170
rect 1665 1215 1770 1245
rect 1665 1170 1695 1215
rect 1740 1170 1770 1215
rect 1665 1140 1770 1170
rect 1905 1200 2010 1230
rect 1905 1155 1935 1200
rect 1980 1155 2010 1200
rect 1905 1125 2010 1155
rect 135 1065 180 1095
rect 1710 1065 1755 1095
rect 135 990 180 1020
rect 1500 990 1545 1020
rect 1710 990 1755 1020
rect 1980 990 2025 1020
rect 1500 915 1545 945
rect 1980 915 2025 945
rect 510 675 615 705
rect 1875 675 1920 705
rect 315 285 360 630
rect 510 630 540 675
rect 585 630 615 675
rect 510 600 615 630
rect 420 495 465 525
rect 420 420 465 450
rect 555 480 600 510
rect 315 210 360 240
rect 420 285 465 315
rect 420 210 465 240
rect 555 285 600 435
rect 555 180 600 240
rect 720 480 765 630
rect 930 615 1035 645
rect 930 570 960 615
rect 1005 570 1035 615
rect 930 540 1035 570
rect 720 285 765 435
rect 960 330 1005 540
rect 1080 495 1125 525
rect 720 210 765 240
rect 1080 180 1125 450
rect 1290 420 1395 450
rect 1290 375 1320 420
rect 1365 375 1395 420
rect 1290 345 1395 375
rect 1215 285 1260 315
rect 1215 210 1260 240
rect 1605 285 1650 630
rect 1875 600 1920 630
rect 1605 210 1650 240
rect 1710 270 1755 300
rect 1710 195 1755 225
rect 1875 270 1920 300
rect 1875 195 1920 225
rect 705 135 810 165
rect 705 90 735 135
rect 780 90 810 135
rect 705 60 810 90
rect 1065 150 1170 180
rect 1065 105 1095 150
rect 1140 105 1170 150
rect 1065 75 1170 105
rect 1335 150 1380 180
rect 1335 75 1380 105
rect 1980 150 2025 180
rect 1980 75 2025 105
<< viali >>
rect 270 1245 315 1290
rect 120 1170 165 1215
rect 435 1155 480 1200
rect 1515 1170 1560 1215
rect 1695 1170 1740 1215
rect 1935 1155 1980 1200
rect 135 1020 180 1065
rect 1710 1020 1755 1065
rect 1500 945 1545 990
rect 1980 945 2025 990
rect 315 630 360 675
rect 540 630 585 675
rect 720 630 765 675
rect 420 450 465 495
rect 420 240 465 285
rect 1605 630 1650 675
rect 960 285 1005 330
rect 1080 450 1125 495
rect 1320 375 1365 420
rect 1215 240 1260 285
rect 1875 630 1920 675
rect 1710 225 1755 270
rect 1875 225 1920 270
rect 555 135 600 180
rect 735 90 780 135
rect 1335 105 1380 150
rect 1980 105 2025 150
<< metal1 >>
rect 255 1290 330 1305
rect 255 1245 270 1290
rect 315 1245 330 1290
rect 255 1230 330 1245
rect 105 1215 180 1230
rect 1500 1215 1575 1230
rect 105 1170 120 1215
rect 165 1170 180 1215
rect 105 1155 180 1170
rect 420 1200 495 1215
rect 420 1155 435 1200
rect 480 1155 495 1200
rect 1500 1170 1515 1215
rect 1560 1170 1575 1215
rect 1500 1155 1575 1170
rect 1680 1215 1755 1230
rect 1680 1170 1695 1215
rect 1740 1170 1755 1215
rect 1680 1155 1755 1170
rect 1920 1200 1995 1215
rect 1920 1155 1935 1200
rect 1980 1155 1995 1200
rect 420 1140 495 1155
rect 1920 1140 1995 1155
rect 120 1065 1770 1080
rect 120 1020 135 1065
rect 180 1050 1710 1065
rect 180 1020 195 1050
rect 120 1005 195 1020
rect 1695 1020 1710 1050
rect 1755 1020 1770 1065
rect 1695 1005 1770 1020
rect 1485 990 1560 1005
rect 1485 945 1500 990
rect 1545 960 1560 990
rect 1965 990 2040 1005
rect 1965 960 1980 990
rect 1545 945 1980 960
rect 2025 945 2040 990
rect 1485 930 2040 945
rect 300 675 1935 690
rect 300 630 315 675
rect 360 660 540 675
rect 360 630 375 660
rect 300 615 375 630
rect 525 630 540 660
rect 585 660 720 675
rect 585 630 600 660
rect 525 615 600 630
rect 705 630 720 660
rect 765 660 1605 675
rect 765 630 780 660
rect 705 615 780 630
rect 1590 630 1605 660
rect 1650 660 1875 675
rect 1650 630 1665 660
rect 1590 615 1665 630
rect 1860 630 1875 660
rect 1920 630 1935 675
rect 1860 615 1935 630
rect 405 495 480 510
rect 1065 495 1140 510
rect 405 450 420 495
rect 465 465 1080 495
rect 465 450 480 465
rect 405 435 480 450
rect 1065 450 1080 465
rect 1125 450 1140 495
rect 1065 435 1140 450
rect 1305 420 1380 435
rect 1305 375 1320 420
rect 1365 375 1380 420
rect 1305 360 1380 375
rect 945 330 1020 345
rect 945 300 960 330
rect 405 285 960 300
rect 1005 300 1020 330
rect 1005 285 1275 300
rect 405 240 420 285
rect 465 270 1215 285
rect 465 240 480 270
rect 405 225 480 240
rect 1200 240 1215 270
rect 1260 240 1275 285
rect 1200 225 1275 240
rect 1695 270 1935 285
rect 1695 225 1710 270
rect 1755 255 1875 270
rect 1755 225 1770 255
rect 1695 210 1770 225
rect 1860 225 1875 255
rect 1920 225 1935 270
rect 1860 210 1935 225
rect 540 180 615 195
rect 540 135 555 180
rect 600 150 615 180
rect 1320 150 2040 165
rect 600 135 795 150
rect 540 120 735 135
rect 720 90 735 120
rect 780 90 795 135
rect 1320 105 1335 150
rect 1380 135 1980 150
rect 1380 105 1395 135
rect 1320 90 1395 105
rect 1965 105 1980 135
rect 2025 105 2040 150
rect 1965 90 2040 105
rect 720 75 795 90
<< labels >>
rlabel pdiff 1067 422 1067 422 3 Vdd
flabel pdiff 165 420 165 420 1 FreeSerif 120 0 0 0 #11
flabel poly 195 405 195 405 3 FreeSerif 120 0 0 0 in(2)
flabel poly 270 405 270 405 3 FreeSerif 120 0 0 0 in(1)
flabel poly 375 360 375 360 3 FreeSerif 120 0 0 0 in(0)
flabel poly 480 360 480 360 3 FreeSerif 120 0 0 0 out
flabel pdiff 450 420 450 420 1 FreeSerif 120 0 0 0 Vdd
flabel pdiff 585 420 585 420 1 FreeSerif 120 0 0 0 #17
flabel poly 780 360 780 360 3 FreeSerif 120 0 0 0 #17
flabel pdiff 750 420 750 420 1 FreeSerif 120 0 0 0 out
flabel poly 885 405 885 405 3 FreeSerif 120 0 0 0 GND
flabel poly 885 315 885 315 3 FreeSerif 120 0 0 0 Vdd
flabel pdiff 1110 420 1110 420 1 FreeSerif 120 0 0 0 Vdd
flabel poly 1290 315 1290 315 3 FreeSerif 120 0 0 0 in(6)
flabel poly 1560 405 1560 405 3 FreeSerif 120 0 0 0 in(4)
flabel pdiff 1530 420 1530 420 1 FreeSerif 120 0 0 0 #9
flabel pdiff 1740 420 1740 420 1 FreeSerif 120 0 0 0 #11
flabel poly 1665 360 1665 360 3 FreeSerif 120 0 0 0 in(3)
flabel poly 1935 360 1935 360 3 FreeSerif 120 0 0 0 in(5)
flabel pdiff 2010 420 2010 420 1 FreeSerif 120 0 0 0 #9
flabel pdiff 1905 420 1905 420 1 FreeSerif 120 0 0 0 out
flabel ndiff 1905 75 1905 75 1 FreeSerif 120 0 0 0 #4
flabel ndiff 1740 75 1740 75 1 FreeSerif 120 0 0 0 #4
flabel ndiff 1635 75 1635 75 1 FreeSerif 120 0 0 0 out
flabel ndiff 1365 75 1365 75 1 FreeSerif 120 0 0 0 #5
flabel ndiff 1215 210 1215 210 1 FreeSerif 120 0 0 0 GND
flabel ndiff 750 210 750 210 1 FreeSerif 120 0 0 0 out
flabel ndiff 345 210 345 210 1 FreeSerif 120 0 0 0 out
flabel ndiff 450 210 450 210 1 FreeSerif 120 0 0 0 GND
flabel ndiff 585 210 585 210 1 FreeSerif 120 0 0 0 #17
flabel ndiff 2010 75 2010 75 1 FreeSerif 120 0 0 0 #5
flabel metal1 990 345 990 345 1 FreeSerif 120 0 0 0 GND
port 1 n
flabel metal1 1125 510 1125 510 1 FreeSerif 120 0 0 0 Vdd
port 2 n
flabel metal1 1350 435 1350 435 1 FreeSerif 120 0 0 0 in(6)
port 3 n
flabel metal1 1965 1215 1965 1215 1 FreeSerif 120 0 0 0 in(5)
port 4 n
flabel metal1 1530 1230 1530 1230 1 FreeSerif 120 0 0 0 in(4)
port 5 n
flabel metal1 1725 1230 1725 1230 1 FreeSerif 120 0 0 0 in(3)
port 6 n
flabel metal1 135 1230 135 1230 1 FreeSerif 120 0 0 0 in(2)
port 7 n
flabel metal1 285 1305 285 1305 1 FreeSerif 120 0 0 0 in(1)
port 8 n
flabel metal1 570 690 570 690 1 FreeSerif 120 0 0 0 out
port 9 n
flabel metal1 465 1215 465 1215 1 FreeSerif 120 0 0 0 in(0)
port 10 n
<< end >>
