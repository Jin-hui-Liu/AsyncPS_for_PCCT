magic
tech sky130A
magscale 1 2
timestamp 1753210778
<< nwell >>
rect 75 555 435 750
rect 75 315 583 555
rect 1125 495 1380 750
rect 1125 315 1755 495
<< nmos >>
rect 300 150 330 240
rect 405 150 465 240
rect 705 150 1035 240
rect 1140 90 1170 240
rect 1245 90 1275 240
rect 1350 150 1380 240
<< pmos >>
rect 195 360 225 705
rect 300 360 330 705
rect 405 360 465 510
rect 1245 360 1275 705
rect 1350 360 1380 450
rect 1425 360 1635 450
<< ndiff >>
rect 225 225 300 240
rect 225 180 240 225
rect 285 180 300 225
rect 225 150 300 180
rect 330 210 405 240
rect 330 165 345 210
rect 390 165 405 210
rect 330 150 405 165
rect 465 225 540 240
rect 465 180 480 225
rect 525 180 540 225
rect 465 150 540 180
rect 630 225 705 240
rect 630 180 645 225
rect 690 180 705 225
rect 630 150 705 180
rect 1035 210 1140 240
rect 1035 165 1065 210
rect 1110 165 1140 210
rect 1035 150 1140 165
rect 1080 90 1140 150
rect 1170 90 1245 240
rect 1275 225 1350 240
rect 1275 180 1290 225
rect 1335 180 1350 225
rect 1275 150 1350 180
rect 1380 225 1455 240
rect 1380 180 1395 225
rect 1440 180 1455 225
rect 1380 150 1455 180
rect 1275 90 1335 150
<< pdiff >>
rect 120 660 195 705
rect 120 615 135 660
rect 180 615 195 660
rect 120 360 195 615
rect 225 360 300 705
rect 330 510 390 705
rect 1170 660 1245 705
rect 1170 615 1185 660
rect 1230 615 1245 660
rect 330 435 405 510
rect 330 390 345 435
rect 390 390 405 435
rect 330 360 405 390
rect 465 420 540 510
rect 465 375 480 420
rect 525 375 540 420
rect 465 360 540 375
rect 1170 360 1245 615
rect 1275 450 1335 705
rect 1275 420 1350 450
rect 1275 375 1290 420
rect 1335 375 1350 420
rect 1275 360 1350 375
rect 1380 360 1425 450
rect 1635 435 1710 450
rect 1635 390 1650 435
rect 1695 390 1710 435
rect 1635 360 1710 390
<< ndiffc >>
rect 240 180 285 225
rect 345 165 390 210
rect 480 180 525 225
rect 645 180 690 225
rect 1065 165 1110 210
rect 1290 180 1335 225
rect 1395 180 1440 225
<< pdiffc >>
rect 135 615 180 660
rect 1185 615 1230 660
rect 345 390 390 435
rect 480 375 525 420
rect 1290 375 1335 420
rect 1650 390 1695 435
<< poly >>
rect 120 810 225 840
rect 120 765 150 810
rect 195 765 225 810
rect 120 735 225 765
rect 195 705 225 735
rect 300 810 405 840
rect 300 765 330 810
rect 375 765 405 810
rect 300 735 405 765
rect 1200 810 1305 840
rect 1200 765 1230 810
rect 1275 765 1305 810
rect 1200 735 1305 765
rect 300 705 330 735
rect 1245 705 1275 735
rect 405 615 525 645
rect 405 570 450 615
rect 495 570 525 615
rect 405 540 525 570
rect 405 510 465 540
rect 810 375 915 405
rect 195 330 225 360
rect 300 240 330 360
rect 405 240 465 360
rect 810 330 840 375
rect 885 330 915 375
rect 1350 600 1485 630
rect 1350 555 1410 600
rect 1455 555 1485 600
rect 1350 525 1485 555
rect 1350 450 1380 525
rect 1425 450 1635 480
rect 810 270 915 330
rect 705 240 1035 270
rect 1140 240 1170 270
rect 1245 240 1275 360
rect 1350 240 1380 360
rect 1425 330 1635 360
rect 1485 300 1590 330
rect 1485 255 1515 300
rect 1560 255 1590 300
rect 300 120 330 150
rect 405 120 465 150
rect 705 120 1035 150
rect 1485 225 1590 255
rect 1350 120 1380 150
rect 1140 0 1170 90
rect 1245 60 1275 90
rect 1140 -30 1245 0
rect 1140 -75 1170 -30
rect 1215 -75 1245 -30
rect 1140 -105 1245 -75
<< polycont >>
rect 150 765 195 810
rect 330 765 375 810
rect 1230 765 1275 810
rect 450 570 495 615
rect 840 330 885 375
rect 1410 555 1455 600
rect 1515 255 1560 300
rect 1170 -75 1215 -30
<< locali >>
rect 120 810 225 840
rect 120 765 150 810
rect 195 765 225 810
rect 120 735 225 765
rect 300 810 405 840
rect 300 765 330 810
rect 375 765 405 810
rect 300 735 405 765
rect 1200 810 1305 840
rect 1200 765 1230 810
rect 1275 765 1305 810
rect 1200 735 1305 765
rect 135 660 180 690
rect 1185 660 1230 690
rect 135 585 180 615
rect 420 615 525 645
rect 420 570 450 615
rect 495 570 525 615
rect 1185 585 1230 615
rect 1380 600 1485 630
rect 420 540 525 570
rect 1380 555 1410 600
rect 1455 555 1485 600
rect 240 225 285 525
rect 1380 525 1485 555
rect 345 435 390 465
rect 345 360 390 390
rect 480 420 525 450
rect 1290 420 1335 510
rect 240 150 285 180
rect 345 210 390 240
rect 345 120 390 165
rect 480 225 525 375
rect 810 375 915 405
rect 810 330 840 375
rect 885 330 915 375
rect 810 300 915 330
rect 480 150 525 180
rect 645 225 690 255
rect 645 150 690 180
rect 1065 210 1110 240
rect 1065 75 1110 165
rect 1290 225 1335 375
rect 1650 435 1695 465
rect 1650 360 1695 390
rect 1485 300 1590 330
rect 1485 255 1515 300
rect 1560 255 1590 300
rect 1290 150 1335 180
rect 1395 225 1440 255
rect 1485 225 1590 255
rect 1395 150 1440 180
rect 1140 -30 1245 0
rect 1140 -75 1170 -30
rect 1215 -75 1245 -30
rect 1140 -105 1245 -75
<< viali >>
rect 150 765 195 810
rect 330 765 375 810
rect 1230 765 1275 810
rect 135 615 180 660
rect 450 570 495 615
rect 1185 615 1230 660
rect 240 525 285 570
rect 1410 555 1455 600
rect 1290 510 1335 555
rect 345 390 390 435
rect 480 450 525 495
rect 840 330 885 375
rect 645 180 690 225
rect 345 75 390 120
rect 1650 390 1695 435
rect 1515 255 1560 300
rect 1395 180 1440 225
rect 1065 30 1110 75
rect 1170 -75 1215 -30
<< metal1 >>
rect 135 810 210 825
rect 135 765 150 810
rect 195 765 210 810
rect 135 750 210 765
rect 315 810 390 825
rect 315 765 330 810
rect 375 765 390 810
rect 315 750 390 765
rect 1215 810 1290 825
rect 1215 765 1230 810
rect 1275 765 1290 810
rect 1215 750 1290 765
rect 120 660 1245 690
rect 120 615 135 660
rect 180 615 195 660
rect 120 600 195 615
rect 435 615 510 630
rect 435 585 450 615
rect 225 570 450 585
rect 495 570 510 615
rect 1170 615 1185 660
rect 1230 615 1245 660
rect 1170 600 1245 615
rect 1395 600 1470 615
rect 225 525 240 570
rect 285 555 1350 570
rect 285 525 300 555
rect 435 540 1290 555
rect 225 510 300 525
rect 1275 510 1290 540
rect 1335 510 1350 555
rect 465 495 540 510
rect 1275 495 1350 510
rect 1395 555 1410 600
rect 1455 555 1470 600
rect 1395 540 1470 555
rect 465 450 480 495
rect 525 465 540 495
rect 1395 465 1425 540
rect 525 450 1425 465
rect 330 435 405 450
rect 465 435 1425 450
rect 1635 435 1710 450
rect 330 390 345 435
rect 390 405 405 435
rect 1635 405 1650 435
rect 390 390 1650 405
rect 1695 390 1710 435
rect 330 375 1710 390
rect 825 330 840 375
rect 885 330 900 375
rect 825 315 900 330
rect 1500 300 1575 315
rect 1500 255 1515 300
rect 1560 255 1575 300
rect 1500 240 1575 255
rect 630 225 705 240
rect 630 180 645 225
rect 690 210 705 225
rect 1380 225 1455 240
rect 1380 210 1395 225
rect 690 180 1395 210
rect 1440 180 1455 225
rect 630 165 705 180
rect 1380 165 1455 180
rect 330 120 405 135
rect 330 75 345 120
rect 390 90 405 120
rect 1500 90 1530 240
rect 390 75 1530 90
rect 330 60 1065 75
rect 1050 30 1065 60
rect 1110 60 1530 75
rect 1110 30 1125 60
rect 1050 15 1125 30
rect 1155 -30 1230 -15
rect 1155 -75 1170 -30
rect 1215 -75 1230 -30
rect 1155 -90 1230 -75
<< labels >>
flabel poly 1245 285 1245 285 3 FreeSerif 120 0 0 0 in(2)
flabel poly 1350 285 1350 285 3 FreeSerif 120 0 0 0 #10
flabel poly 720 255 720 255 3 FreeSerif 120 0 0 0 Vdd
rlabel poly 197 332 197 332 3 in(1)
rlabel poly 1427 332 1427 332 3 GND
flabel poly 300 330 300 330 3 FreeSerif 120 0 0 0 in(0)
flabel poly 405 315 405 315 3 FreeSerif 120 0 0 0 out
flabel pdiff 120 375 120 375 3 FreeSerif 120 0 0 0 #7
flabel pdiff 345 375 345 375 3 FreeSerif 120 0 0 0 Vdd
flabel pdiff 480 375 480 375 3 FreeSerif 120 0 0 0 #10
flabel pdiff 1185 375 1185 375 3 FreeSerif 120 0 0 0 #7
flabel pdiff 1290 375 1290 375 3 FreeSerif 120 0 0 0 out
flabel pdiff 1650 375 1650 375 3 FreeSerif 120 0 0 0 Vdd
flabel poly 1440 330 1440 330 1 FreeSerif 120 0 0 0 GND
flabel ndiff 1395 165 1395 165 3 FreeSerif 120 0 0 0 #12
flabel ndiff 1290 105 1290 105 3 FreeSerif 120 0 0 0 out
flabel poly 1140 255 1140 255 3 FreeSerif 120 0 0 0 in(3)
flabel ndiff 1050 165 1050 165 3 FreeSerif 120 0 0 0 GND
flabel ndiff 645 165 645 165 3 FreeSerif 120 0 0 0 #12
flabel ndiff 480 165 480 165 3 FreeSerif 120 0 0 0 #10
flabel ndiff 240 165 240 165 3 FreeSerif 120 0 0 0 out
flabel poly 195 345 195 345 3 FreeSerif 120 0 0 0 in(1)
flabel ndiff 345 180 345 180 3 FreeSerif 120 0 0 0 GND
flabel metal1 165 825 165 825 1 FreeSerif 120 0 0 0 in(1)
port 5 n
flabel metal1 360 825 360 825 1 FreeSerif 120 0 0 0 in(0)
port 7 n
flabel metal1 1230 -60 1230 -60 3 FreeSerif 120 0 0 0 in(3)
port 3 e
flabel metal1 1245 825 1245 825 1 FreeSerif 120 0 0 0 in(2)
port 4 n
flabel metal1 1575 270 1575 270 3 FreeSerif 120 0 0 0 GND
port 1 e
flabel metal1 510 600 510 600 3 FreeSerif 120 0 0 0 out
port 6 e
flabel metal1 855 405 855 405 1 FreeSerif 120 0 0 0 Vdd
port 2 n
<< end >>
