magic
tech sky130A
magscale 1 2
timestamp 1753015928
<< checkpaint >>
rect -1140 2205 2400 2280
rect -1140 2175 2985 2205
rect -1140 -1200 3060 2175
rect -1065 -1230 2985 -1200
<< nmos >>
rect 195 60 225 360
rect 300 60 330 360
rect 405 270 435 360
rect 510 270 570 360
rect 915 270 945 360
rect 990 270 1320 360
rect 1425 60 1455 360
rect 1695 60 1725 360
<< pmos >>
rect 300 465 330 915
rect 405 465 435 915
rect 510 465 570 615
rect 810 465 840 915
rect 915 465 945 555
rect 990 465 1200 555
rect 1695 465 1725 915
<< ndiff >>
rect 120 60 195 360
rect 225 60 300 360
rect 330 270 405 360
rect 435 270 510 360
rect 570 270 645 360
rect 840 270 915 360
rect 945 270 990 360
rect 1320 270 1425 360
rect 330 60 390 270
rect 1365 60 1425 270
rect 1455 60 1530 360
rect 1620 60 1695 360
rect 1725 60 1800 360
<< pdiff >>
rect 225 465 300 915
rect 330 465 405 915
rect 435 615 495 915
rect 435 465 510 615
rect 570 465 645 615
rect 735 465 810 915
rect 840 555 900 915
rect 840 465 915 555
rect 945 465 990 555
rect 1200 465 1275 555
rect 1620 465 1695 915
rect 1725 465 1800 915
<< poly >>
rect 300 915 330 945
rect 405 915 435 945
rect 810 915 840 945
rect 1695 915 1725 945
rect 510 615 570 645
rect 915 555 945 585
rect 990 555 1200 585
rect 300 435 330 465
rect 405 435 435 465
rect 510 435 570 465
rect 810 435 840 465
rect 915 435 945 465
rect 990 435 1200 465
rect 1695 435 1725 465
rect 195 360 225 390
rect 300 360 330 390
rect 405 360 435 390
rect 510 360 570 390
rect 915 360 945 390
rect 990 360 1320 390
rect 1425 360 1455 390
rect 1695 360 1725 390
rect 405 240 435 270
rect 510 240 570 270
rect 915 240 945 270
rect 990 240 1320 270
rect 195 30 225 60
rect 300 30 330 60
rect 1425 30 1455 60
rect 1695 30 1725 60
<< metal1 >>
rect 120 960 180 1020
rect 240 960 300 1020
rect 360 960 420 1020
rect 480 960 540 1020
rect 600 960 660 1020
rect 720 960 780 1020
rect 840 960 900 1020
rect 960 960 1020 1020
rect 1080 960 1140 1020
rect 120 60 180 120
<< labels >>
rlabel ndiff 572 272 572 272 3 #16
rlabel pdiff 572 467 572 467 3 #16
rlabel poly 512 362 512 362 3 out
rlabel poly 512 437 512 437 3 out
rlabel ndiff 437 272 437 272 3 GND
rlabel poly 407 362 407 362 3 in(0)
rlabel poly 407 437 407 437 3 in(0)
rlabel pdiff 437 467 437 467 3 Vdd
rlabel ndiff 332 62 332 62 3 out
rlabel poly 302 362 302 362 3 in(6)
rlabel poly 302 437 302 437 3 in(1)
rlabel pdiff 227 467 227 467 3 #12
rlabel poly 197 362 197 362 3 in(5)
rlabel ndiff 122 62 122 62 3 #5
rlabel poly 1427 362 1427 362 3 in(4)
rlabel pdiff 1202 467 1202 467 3 Vdd
rlabel ndiff 1457 62 1457 62 3 #6
rlabel ndiff 1322 272 1322 272 3 GND
rlabel poly 992 362 992 362 3 Vdd
rlabel poly 992 437 992 437 3 GND
rlabel poly 917 362 917 362 3 #16
rlabel poly 917 437 917 437 3 #16
rlabel ndiff 842 272 842 272 3 out
rlabel pdiff 842 467 842 467 3 out
rlabel poly 812 437 812 437 3 in(3)
rlabel pdiff 737 467 737 467 3 #11
rlabel ndiff 1727 62 1727 62 3 #6
rlabel pdiff 1727 467 1727 467 3 #11
rlabel poly 1697 362 1697 362 3 in(2)
rlabel poly 1697 437 1697 437 3 in(2)
rlabel ndiff 1622 62 1622 62 3 #5
rlabel pdiff 1622 467 1622 467 3 #12
rlabel metal1 1082 962 1082 962 3 GND
port 1 e
rlabel metal1 962 962 962 962 3 Vdd
port 2 e
rlabel metal1 842 962 842 962 3 in(6)
port 3 e
rlabel metal1 722 962 722 962 3 in(5)
port 4 e
rlabel metal1 602 962 602 962 3 in(4)
port 5 e
rlabel metal1 482 962 482 962 3 in(3)
port 6 e
rlabel metal1 362 962 362 962 3 in(2)
port 7 e
rlabel metal1 242 962 242 962 3 in(1)
port 8 e
rlabel metal1 122 62 122 62 3 out
rlabel metal1 122 962 122 962 3 in(0)
port 9 e
<< end >>
