magic
tech sky130A
magscale 1 2
timestamp 1753015927
<< checkpaint >>
rect -1140 2265 2400 2340
rect -1140 2235 2985 2265
rect -1140 -1185 3060 2235
rect -1140 -1200 2985 -1185
rect -960 -1215 2985 -1200
<< nmos >>
rect 300 75 330 300
rect 405 210 435 300
rect 510 210 570 300
rect 915 210 945 300
rect 990 210 1320 300
rect 1425 75 1455 300
rect 1695 75 1725 300
<< pmos >>
rect 195 405 225 975
rect 300 405 330 975
rect 405 405 435 975
rect 510 405 570 555
rect 810 405 840 975
rect 915 405 945 495
rect 990 405 1200 495
rect 1695 405 1725 975
<< ndiff >>
rect 225 75 300 300
rect 330 210 405 300
rect 435 210 510 300
rect 570 210 645 300
rect 840 210 915 300
rect 945 210 990 300
rect 1320 210 1425 300
rect 330 75 390 210
rect 1365 75 1425 210
rect 1455 75 1530 300
rect 1620 75 1695 300
rect 1725 75 1800 300
<< pdiff >>
rect 120 405 195 975
rect 225 405 300 975
rect 330 405 405 975
rect 435 555 495 975
rect 435 405 510 555
rect 570 405 645 555
rect 735 405 810 975
rect 840 495 900 975
rect 840 405 915 495
rect 945 405 990 495
rect 1200 405 1275 495
rect 1620 405 1695 975
rect 1725 405 1800 975
<< poly >>
rect 195 975 225 1005
rect 300 975 330 1005
rect 405 975 435 1005
rect 810 975 840 1005
rect 1695 975 1725 1005
rect 510 555 570 585
rect 915 495 945 525
rect 990 495 1200 525
rect 195 375 225 405
rect 300 375 330 405
rect 405 375 435 405
rect 510 375 570 405
rect 810 375 840 405
rect 915 375 945 405
rect 990 375 1200 405
rect 1695 375 1725 405
rect 300 300 330 330
rect 405 300 435 330
rect 510 300 570 330
rect 915 300 945 330
rect 990 300 1320 330
rect 1425 300 1455 330
rect 1695 300 1725 330
rect 405 180 435 210
rect 510 180 570 210
rect 915 180 945 210
rect 990 180 1320 210
rect 300 45 330 75
rect 1425 45 1455 75
rect 1695 45 1725 75
<< metal1 >>
rect 120 1020 180 1080
rect 240 1020 300 1080
rect 360 1020 420 1080
rect 480 1020 540 1080
rect 600 1020 660 1080
rect 720 1020 780 1080
rect 840 1020 900 1080
rect 960 1020 1020 1080
rect 1080 1020 1140 1080
rect 120 60 180 120
<< labels >>
rlabel ndiff 572 212 572 212 3 #16
rlabel pdiff 572 407 572 407 3 #16
rlabel poly 512 302 512 302 3 out
rlabel ndiff 437 212 437 212 3 GND
rlabel poly 512 377 512 377 3 out
rlabel poly 407 302 407 302 3 in(0)
rlabel pdiff 437 407 437 407 3 Vdd
rlabel poly 407 377 407 377 3 in(0)
rlabel ndiff 332 77 332 77 3 out
rlabel poly 302 302 302 302 3 in(6)
rlabel poly 302 377 302 377 3 in(1)
rlabel ndiff 227 77 227 77 3 #4
rlabel poly 197 377 197 377 3 in(2)
rlabel pdiff 122 407 122 407 3 #10
rlabel poly 1427 302 1427 302 3 in(5)
rlabel pdiff 1202 407 1202 407 3 Vdd
rlabel ndiff 1457 77 1457 77 3 #5
rlabel ndiff 1322 212 1322 212 3 GND
rlabel poly 992 302 992 302 3 Vdd
rlabel poly 992 377 992 377 3 GND
rlabel poly 917 302 917 302 3 #16
rlabel poly 917 377 917 377 3 #16
rlabel ndiff 842 212 842 212 3 out
rlabel pdiff 842 407 842 407 3 out
rlabel poly 812 377 812 377 3 in(4)
rlabel pdiff 737 407 737 407 3 #9
rlabel ndiff 1727 77 1727 77 3 #5
rlabel pdiff 1727 407 1727 407 3 #9
rlabel poly 1697 302 1697 302 3 in(3)
rlabel poly 1697 377 1697 377 3 in(3)
rlabel ndiff 1622 77 1622 77 3 #4
rlabel pdiff 1622 407 1622 407 3 #10
rlabel metal1 1082 1022 1082 1022 3 GND
port 1 e
rlabel metal1 962 1022 962 1022 3 Vdd
port 2 e
rlabel metal1 842 1022 842 1022 3 in(6)
port 3 e
rlabel metal1 722 1022 722 1022 3 in(5)
port 4 e
rlabel metal1 602 1022 602 1022 3 in(4)
port 5 e
rlabel metal1 482 1022 482 1022 3 in(3)
port 6 e
rlabel metal1 362 1022 362 1022 3 in(2)
port 7 e
rlabel metal1 242 1022 242 1022 3 in(1)
port 8 e
rlabel metal1 122 62 122 62 3 out
port 9 e
rlabel metal1 122 1022 122 1022 3 in(0)
port 10 e
<< end >>
