magic
tech sky130A
magscale 1 2
timestamp 1753291491
<< nwell >>
rect 360 975 750 1110
rect 360 825 1530 975
rect 360 765 2040 825
rect 225 615 2040 765
rect 75 495 2040 615
rect 75 315 2415 495
<< nmos >>
rect 720 150 1050 240
rect 1155 90 1185 240
rect 1260 90 1290 240
rect 1395 150 1425 240
rect 1500 150 1560 240
rect 1800 90 1830 240
rect 1905 90 1935 240
rect 2010 150 2040 240
<< pmos >>
rect 195 360 225 570
rect 330 360 360 720
rect 465 360 495 1065
rect 540 360 570 1065
rect 615 360 645 1065
rect 720 360 750 930
rect 1155 360 1185 930
rect 1260 360 1290 645
rect 1395 360 1425 930
rect 1500 360 1560 510
rect 1905 360 1935 780
rect 2010 360 2040 450
rect 2085 360 2295 450
<< ndiff >>
rect 645 210 720 240
rect 645 165 660 210
rect 705 165 720 210
rect 645 150 720 165
rect 1050 210 1155 240
rect 1050 165 1080 210
rect 1125 165 1155 210
rect 1050 150 1155 165
rect 1095 90 1155 150
rect 1185 90 1260 240
rect 1290 225 1395 240
rect 1290 180 1335 225
rect 1380 180 1395 225
rect 1290 150 1395 180
rect 1425 210 1500 240
rect 1425 165 1440 210
rect 1485 165 1500 210
rect 1425 150 1500 165
rect 1560 225 1635 240
rect 1560 180 1575 225
rect 1620 180 1635 225
rect 1560 150 1635 180
rect 1725 150 1800 240
rect 1290 90 1350 150
rect 1725 105 1740 150
rect 1785 105 1800 150
rect 1725 90 1800 105
rect 1830 90 1905 240
rect 1935 225 2010 240
rect 1935 180 1950 225
rect 1995 180 2010 225
rect 1935 150 2010 180
rect 2040 210 2115 240
rect 2040 165 2055 210
rect 2100 165 2115 210
rect 2040 150 2115 165
rect 1935 90 1995 150
<< pdiff >>
rect 405 720 465 1065
rect 270 570 330 720
rect 120 435 195 570
rect 120 390 135 435
rect 180 390 195 435
rect 120 360 195 390
rect 225 510 330 570
rect 225 465 255 510
rect 300 465 330 510
rect 225 360 330 465
rect 360 360 465 720
rect 495 360 540 1065
rect 570 360 615 1065
rect 645 930 705 1065
rect 645 720 720 930
rect 645 675 660 720
rect 705 675 720 720
rect 645 360 720 675
rect 750 360 1155 930
rect 1185 645 1245 930
rect 1335 645 1395 930
rect 1185 360 1260 645
rect 1290 615 1395 645
rect 1290 570 1305 615
rect 1350 570 1395 615
rect 1290 360 1395 570
rect 1425 510 1485 930
rect 1425 495 1500 510
rect 1425 450 1440 495
rect 1485 450 1500 495
rect 1425 360 1500 450
rect 1560 420 1635 510
rect 1560 375 1575 420
rect 1620 375 1635 420
rect 1560 360 1635 375
rect 1830 435 1905 780
rect 1830 390 1845 435
rect 1890 390 1905 435
rect 1830 360 1905 390
rect 1935 450 1995 780
rect 1935 420 2010 450
rect 1935 375 1950 420
rect 1995 375 2010 420
rect 1935 360 2010 375
rect 2040 360 2085 450
rect 2295 420 2370 450
rect 2295 375 2310 420
rect 2355 375 2370 420
rect 2295 360 2370 375
<< ndiffc >>
rect 660 165 705 210
rect 1080 165 1125 210
rect 1335 180 1380 225
rect 1440 165 1485 210
rect 1575 180 1620 225
rect 1740 105 1785 150
rect 1950 180 1995 225
rect 2055 165 2100 210
<< pdiffc >>
rect 135 390 180 435
rect 255 465 300 510
rect 660 675 705 720
rect 1305 570 1350 615
rect 1440 450 1485 495
rect 1575 375 1620 420
rect 1845 390 1890 435
rect 1950 375 1995 420
rect 2310 375 2355 420
<< poly >>
rect 465 1260 570 1290
rect 465 1215 495 1260
rect 540 1215 570 1260
rect 315 1170 420 1200
rect 465 1185 570 1215
rect 315 1125 345 1170
rect 390 1125 420 1170
rect 315 1095 495 1125
rect 465 1065 495 1095
rect 540 1065 570 1185
rect 615 1260 720 1290
rect 615 1215 645 1260
rect 690 1215 720 1260
rect 615 1185 720 1215
rect 615 1065 645 1185
rect 270 825 375 855
rect 270 780 300 825
rect 345 780 375 825
rect 270 750 375 780
rect 330 720 360 750
rect 135 675 240 705
rect 135 630 165 675
rect 210 630 240 675
rect 135 600 240 630
rect 195 570 225 600
rect 720 1035 855 1065
rect 720 990 780 1035
rect 825 990 855 1035
rect 720 960 855 990
rect 1050 1035 1185 1065
rect 1050 990 1080 1035
rect 1125 990 1185 1035
rect 1050 960 1185 990
rect 1230 1035 1335 1065
rect 1230 990 1260 1035
rect 1305 990 1335 1035
rect 1230 960 1335 990
rect 1395 1035 1530 1065
rect 1395 990 1455 1035
rect 1500 990 1530 1035
rect 1395 960 1530 990
rect 720 930 750 960
rect 1155 930 1185 960
rect 1260 645 1290 960
rect 1395 930 1425 960
rect 1875 885 1980 915
rect 1875 840 1905 885
rect 1950 840 1980 885
rect 1875 810 1980 840
rect 1905 780 1935 810
rect 1530 675 1635 705
rect 1530 630 1560 675
rect 1605 630 1635 675
rect 1530 600 1635 630
rect 1530 570 1575 600
rect 1500 510 1560 570
rect 2040 600 2145 630
rect 2040 555 2070 600
rect 2115 555 2145 600
rect 2010 525 2145 555
rect 2010 450 2040 525
rect 2085 450 2295 480
rect 195 330 225 360
rect 330 330 360 360
rect 465 330 495 360
rect 540 330 570 360
rect 615 330 645 360
rect 720 330 750 360
rect 1155 330 1185 360
rect 720 240 1050 270
rect 1155 240 1185 270
rect 1260 240 1290 360
rect 1395 240 1425 360
rect 1500 240 1560 360
rect 1800 240 1830 270
rect 1905 240 1935 360
rect 2010 240 2040 360
rect 2085 330 2295 360
rect 2145 300 2250 330
rect 2145 255 2175 300
rect 2220 255 2250 300
rect 720 120 1050 150
rect 825 90 930 120
rect 1395 120 1425 150
rect 1500 120 1560 150
rect 2145 225 2250 255
rect 2010 120 2040 150
rect 825 45 855 90
rect 900 45 930 90
rect 1155 45 1185 90
rect 1260 60 1290 90
rect 825 15 930 45
rect 1110 15 1215 45
rect 1110 -30 1140 15
rect 1185 -30 1215 15
rect 1110 -60 1215 -30
rect 1800 0 1830 90
rect 1905 60 1935 90
rect 1800 -30 1905 0
rect 1800 -75 1830 -30
rect 1875 -75 1905 -30
rect 1800 -105 1905 -75
<< polycont >>
rect 495 1215 540 1260
rect 345 1125 390 1170
rect 645 1215 690 1260
rect 300 780 345 825
rect 165 630 210 675
rect 780 990 825 1035
rect 1080 990 1125 1035
rect 1260 990 1305 1035
rect 1455 990 1500 1035
rect 1905 840 1950 885
rect 1560 630 1605 675
rect 2070 555 2115 600
rect 2175 255 2220 300
rect 855 45 900 90
rect 1140 -30 1185 15
rect 1830 -75 1875 -30
<< locali >>
rect 465 1260 570 1290
rect 465 1215 495 1260
rect 540 1215 570 1260
rect 315 1170 420 1200
rect 465 1185 570 1215
rect 615 1260 720 1290
rect 615 1215 645 1260
rect 690 1215 720 1260
rect 615 1185 720 1215
rect 315 1125 345 1170
rect 390 1125 420 1170
rect 315 1095 420 1125
rect 750 1035 855 1065
rect 750 990 780 1035
rect 825 990 855 1035
rect 750 960 855 990
rect 1050 1035 1155 1065
rect 1050 990 1080 1035
rect 1125 990 1155 1035
rect 1050 960 1155 990
rect 1230 1035 1335 1065
rect 1230 990 1260 1035
rect 1305 990 1335 1035
rect 1230 960 1335 990
rect 1425 1035 1530 1065
rect 1425 990 1455 1035
rect 1500 990 1530 1035
rect 1425 960 1530 990
rect 1875 885 1980 915
rect 270 825 375 855
rect 270 780 300 825
rect 345 780 375 825
rect 1875 840 1905 885
rect 1950 840 1980 885
rect 1875 810 1980 840
rect 270 750 375 780
rect 660 720 705 750
rect 135 675 240 705
rect 135 630 165 675
rect 210 630 240 675
rect 660 645 705 675
rect 135 600 240 630
rect 255 510 300 540
rect 135 435 180 465
rect 255 435 300 465
rect 135 360 180 390
rect 660 210 705 240
rect 660 135 705 165
rect 855 120 900 735
rect 1305 615 1350 645
rect 1305 540 1350 570
rect 1440 495 1485 765
rect 1530 675 1635 705
rect 1530 630 1560 675
rect 1605 630 1635 675
rect 1530 600 1635 630
rect 1080 210 1125 240
rect 1080 135 1125 165
rect 1335 225 1380 450
rect 1440 420 1485 450
rect 1575 420 1620 510
rect 1335 150 1380 180
rect 1440 210 1485 240
rect 825 90 930 120
rect 1440 135 1485 165
rect 1575 225 1620 375
rect 1845 435 1890 465
rect 1845 360 1890 390
rect 1950 420 1995 615
rect 2040 600 2145 630
rect 2040 555 2070 600
rect 2115 555 2145 600
rect 2040 525 2145 555
rect 1950 225 1995 375
rect 2310 420 2355 450
rect 2310 345 2355 375
rect 2145 300 2250 330
rect 2145 255 2175 300
rect 2220 255 2250 300
rect 1575 150 1620 180
rect 1740 150 1785 180
rect 1950 150 1995 180
rect 2055 210 2100 240
rect 2145 225 2250 255
rect 2055 135 2100 165
rect 1740 90 1785 105
rect 825 45 855 90
rect 900 45 930 90
rect 825 15 930 45
rect 1110 15 1215 45
rect 1110 -30 1140 15
rect 1185 -30 1215 15
rect 1110 -60 1215 -30
rect 1800 -30 1905 0
rect 1800 -75 1830 -30
rect 1875 -75 1905 -30
rect 1800 -105 1905 -75
<< viali >>
rect 495 1215 540 1260
rect 645 1215 690 1260
rect 345 1125 390 1170
rect 780 990 825 1035
rect 1080 990 1125 1035
rect 1260 990 1305 1035
rect 1455 990 1500 1035
rect 300 780 345 825
rect 1905 840 1950 885
rect 165 630 210 675
rect 660 675 705 720
rect 855 735 900 780
rect 255 465 300 510
rect 135 390 180 435
rect 660 165 705 210
rect 1305 570 1350 615
rect 1560 630 1605 675
rect 1950 615 1995 660
rect 1335 450 1380 495
rect 1575 510 1620 555
rect 1080 90 1125 135
rect 1845 390 1890 435
rect 2070 555 2115 600
rect 2310 375 2355 420
rect 2175 255 2220 300
rect 2055 165 2100 210
rect 1440 90 1485 135
rect 1740 45 1785 90
rect 1140 -30 1185 15
rect 1830 -75 1875 -30
<< metal1 >>
rect 480 1260 555 1275
rect 480 1215 495 1260
rect 540 1215 555 1260
rect 480 1200 555 1215
rect 630 1260 705 1275
rect 630 1215 645 1260
rect 690 1215 705 1260
rect 630 1200 705 1215
rect 330 1170 405 1185
rect 330 1125 345 1170
rect 390 1140 405 1170
rect 390 1125 1920 1140
rect 330 1110 1920 1125
rect 1290 1050 1320 1110
rect 765 1035 840 1050
rect 765 990 780 1035
rect 825 990 840 1035
rect 765 975 840 990
rect 1065 1035 1140 1050
rect 1065 990 1080 1035
rect 1125 990 1140 1035
rect 1065 975 1140 990
rect 1245 1035 1320 1050
rect 1245 990 1260 1035
rect 1305 990 1320 1035
rect 1245 975 1320 990
rect 1440 1035 1515 1050
rect 1440 990 1455 1035
rect 1500 990 1515 1035
rect 1440 975 1515 990
rect 1890 900 1920 1110
rect 1890 885 1965 900
rect 1890 840 1905 885
rect 1950 840 1965 885
rect 285 825 360 840
rect 1890 825 1965 840
rect 285 780 300 825
rect 345 780 360 825
rect 285 765 360 780
rect 840 780 915 795
rect 840 735 855 780
rect 900 765 915 780
rect 900 735 2355 765
rect 645 720 720 735
rect 840 720 915 735
rect 150 675 225 690
rect 150 630 165 675
rect 210 630 225 675
rect 645 675 660 720
rect 705 690 720 720
rect 705 675 1620 690
rect 645 660 1560 675
rect 150 615 225 630
rect 285 615 1365 630
rect 285 600 1305 615
rect 285 525 315 600
rect 1290 570 1305 600
rect 1350 570 1365 615
rect 1290 555 1365 570
rect 1290 540 1320 555
rect 240 510 315 525
rect 1440 510 1470 660
rect 1545 630 1560 660
rect 1605 645 1620 675
rect 1935 660 2010 675
rect 1935 645 1950 660
rect 1605 630 1950 645
rect 1545 615 1950 630
rect 1995 615 2010 660
rect 1935 600 2010 615
rect 2055 600 2130 615
rect 2055 570 2070 600
rect 240 465 255 510
rect 300 465 315 510
rect 240 450 315 465
rect 1320 495 1470 510
rect 1560 555 2070 570
rect 2115 555 2130 600
rect 1560 510 1575 555
rect 1620 540 2130 555
rect 1620 510 1635 540
rect 1560 495 1635 510
rect 1320 450 1335 495
rect 1380 480 1470 495
rect 1380 450 1395 480
rect 120 435 195 450
rect 1320 435 1395 450
rect 1830 435 1905 450
rect 2325 435 2355 735
rect 120 390 135 435
rect 180 405 195 435
rect 1830 405 1845 435
rect 180 390 1845 405
rect 1890 390 1905 435
rect 120 375 1905 390
rect 2295 420 2370 435
rect 2295 375 2310 420
rect 2355 375 2370 420
rect 2295 360 2370 375
rect 2160 300 2235 315
rect 2160 255 2175 300
rect 2220 255 2235 300
rect 2160 240 2235 255
rect 645 210 720 225
rect 2040 210 2115 225
rect 645 165 660 210
rect 705 180 2055 210
rect 705 165 720 180
rect 645 150 720 165
rect 2040 165 2055 180
rect 2100 165 2115 210
rect 2040 150 2115 165
rect 1065 135 1140 150
rect 1065 90 1080 135
rect 1125 105 1140 135
rect 1425 135 1500 150
rect 1425 105 1440 135
rect 1125 90 1440 105
rect 1485 105 1500 135
rect 2205 105 2235 240
rect 1485 90 2235 105
rect 1065 75 1740 90
rect 1725 45 1740 75
rect 1785 75 2235 90
rect 1785 45 1800 75
rect 1725 30 1800 45
rect 1125 15 1200 30
rect 1125 -30 1140 15
rect 1185 -30 1200 15
rect 1125 -45 1200 -30
rect 1815 -30 1890 -15
rect 1815 -75 1830 -30
rect 1875 -75 1890 -30
rect 1815 -90 1890 -75
<< labels >>
flabel poly 735 255 735 255 1 FreeSerif 120 0 0 0 Vdd
flabel ndiff 645 165 645 165 3 FreeSerif 120 0 0 0 #24
flabel ndiff 1095 120 1095 120 3 FreeSerif 120 0 0 0 GND
flabel poly 1155 255 1155 255 3 FreeSerif 120 0 0 0 in(8)
flabel poly 1155 345 1155 345 3 FreeSerif 120 0 0 0 in(6)
flabel ndiff 1350 120 1350 120 7 FreeSerif 120 0 0 0 out
flabel ndiff 1620 150 1620 150 1 FreeSerif 120 0 0 0 #22
flabel ndiff 1485 150 1485 150 1 FreeSerif 120 0 0 0 GND
flabel ndiff 1755 90 1755 90 1 FreeSerif 120 0 0 0 GND
flabel ndiff 1980 90 1980 90 1 FreeSerif 120 0 0 0 out
flabel ndiff 2100 150 2100 150 1 FreeSerif 120 0 0 0 #24
flabel pdiff 2355 360 2355 360 1 FreeSerif 120 0 0 0 Vdd
flabel poly 2115 330 2115 330 1 FreeSerif 120 0 0 0 GND
flabel poly 2010 285 2010 285 3 FreeSerif 120 0 0 0 #22
flabel poly 1905 285 1905 285 3 FreeSerif 120 0 0 0 in(2)
flabel pdiff 1980 360 1980 360 1 FreeSerif 120 0 0 0 out
flabel pdiff 1875 360 1875 360 1 FreeSerif 120 0 0 0 #10
flabel poly 1800 255 1800 255 1 FreeSerif 120 0 0 0 in(9)
flabel poly 1260 285 1260 285 3 FreeSerif 120 0 0 0 in(2)
flabel poly 1395 285 1395 285 3 FreeSerif 120 0 0 0 in(0)
flabel poly 1500 285 1500 285 3 FreeSerif 120 0 0 0 out
flabel pdiff 1620 360 1620 360 1 FreeSerif 120 0 0 0 #22
flabel pdiff 1485 360 1485 360 1 FreeSerif 120 0 0 0 Vdd
flabel pdiff 1365 360 1365 360 1 FreeSerif 120 0 0 0 #9
flabel pdiff 690 360 690 360 1 FreeSerif 120 0 0 0 out
flabel pdiff 300 360 300 360 1 FreeSerif 120 0 0 0 #9
flabel pdiff 180 360 180 360 1 FreeSerif 120 0 0 0 #10
flabel poly 465 345 465 345 3 FreeSerif 120 0 0 0 in(2)
flabel poly 540 345 540 345 3 FreeSerif 120 0 0 0 in(4)
flabel poly 615 345 615 345 3 FreeSerif 120 0 0 0 in(5)
flabel poly 720 345 720 345 3 FreeSerif 120 0 0 0 in(7)
flabel poly 195 345 195 345 3 FreeSerif 120 0 0 0 in(1)
flabel poly 330 345 330 345 3 FreeSerif 120 0 0 0 in(3)
flabel metal1 1155 -45 1155 -45 5 FreeSerif 120 0 0 0 in(8)
port 4 s
flabel metal1 180 690 180 690 1 FreeSerif 120 0 0 0 in(1)
port 11 n
flabel metal1 315 840 315 840 1 FreeSerif 120 0 0 0 in(3)
port 9 n
flabel metal1 510 1275 510 1275 1 FreeSerif 120 0 0 0 in(4)
port 8 n
flabel metal1 675 1275 675 1275 1 FreeSerif 120 0 0 0 in(5)
port 7 n
flabel metal1 1845 -90 1845 -90 5 FreeSerif 120 0 0 0 in(9)
port 3 s
flabel metal1 1275 1050 1275 1050 1 FreeSerif 120 0 0 0 in(2)
port 10 n
flabel metal1 1590 690 1590 690 1 FreeSerif 120 0 0 0 out
port 12 n
flabel metal1 2355 435 2355 435 3 FreeSerif 120 0 0 0 Vdd
port 2 e
flabel metal1 810 1050 810 1050 1 FreeSerif 120 0 0 0 in(7)
port 5 n
flabel metal1 1095 1050 1095 1050 1 FreeSerif 120 0 0 0 in(6)
port 6 n
flabel metal1 1500 1050 1500 1050 1 FreeSerif 120 0 0 0 in(0)
port 13 n
<< end >>
