magic
tech sky130A
magscale 1 2
timestamp 1753015925
<< checkpaint >>
rect -1140 2055 2760 2400
rect -1140 2025 3195 2055
rect -1140 1725 3255 2025
rect -1140 1695 3555 1725
rect -1140 -915 3630 1695
rect -1140 -945 3555 -915
rect -1140 -1110 3375 -945
rect -1140 -1140 3300 -1110
rect -1140 -1170 3255 -1140
rect -1140 -1200 3195 -1170
<< nmos >>
rect 720 150 1050 240
rect 1155 90 1185 240
rect 1260 90 1290 240
rect 1395 150 1425 240
rect 1500 150 1560 240
rect 1800 90 1830 240
rect 1905 90 1935 240
rect 2010 150 2040 240
<< pmos >>
rect 195 345 225 555
rect 330 345 360 705
rect 465 345 495 1050
rect 540 345 570 1050
rect 615 345 645 1050
rect 720 345 750 915
rect 1155 345 1185 915
rect 1260 345 1290 630
rect 1395 345 1425 915
rect 1500 345 1560 495
rect 1905 345 1935 765
rect 2010 345 2040 435
rect 2085 345 2295 435
<< ndiff >>
rect 645 150 720 240
rect 1050 150 1155 240
rect 1095 90 1155 150
rect 1185 90 1260 240
rect 1290 150 1395 240
rect 1425 150 1500 240
rect 1560 150 1635 240
rect 1290 90 1350 150
rect 1725 90 1800 240
rect 1830 90 1905 240
rect 1935 150 2010 240
rect 2040 150 2115 240
rect 1935 90 1995 150
<< pdiff >>
rect 405 705 465 1050
rect 270 555 330 705
rect 120 345 195 555
rect 225 345 330 555
rect 360 345 465 705
rect 495 345 540 1050
rect 570 345 615 1050
rect 645 915 705 1050
rect 645 345 720 915
rect 750 345 1155 915
rect 1185 630 1245 915
rect 1335 630 1395 915
rect 1185 345 1260 630
rect 1290 345 1395 630
rect 1425 495 1485 915
rect 1425 345 1500 495
rect 1560 345 1635 495
rect 1830 345 1905 765
rect 1935 435 1995 765
rect 1935 345 2010 435
rect 2040 345 2085 435
rect 2295 345 2370 435
<< poly >>
rect 465 1050 495 1080
rect 540 1050 570 1080
rect 615 1050 645 1080
rect 330 705 360 735
rect 195 555 225 585
rect 720 915 750 945
rect 1155 915 1185 945
rect 1395 915 1425 945
rect 1260 630 1290 660
rect 1905 765 1935 795
rect 1500 495 1560 525
rect 2010 435 2040 465
rect 2085 435 2295 465
rect 195 315 225 345
rect 330 315 360 345
rect 465 315 495 345
rect 540 315 570 345
rect 615 315 645 345
rect 720 315 750 345
rect 1155 315 1185 345
rect 1260 315 1290 345
rect 1395 315 1425 345
rect 1500 315 1560 345
rect 1905 315 1935 345
rect 2010 315 2040 345
rect 2085 315 2295 345
rect 720 240 1050 270
rect 1155 240 1185 270
rect 1260 240 1290 270
rect 1395 240 1425 270
rect 1500 240 1560 270
rect 1800 240 1830 270
rect 1905 240 1935 270
rect 2010 240 2040 270
rect 720 120 1050 150
rect 1395 120 1425 150
rect 1500 120 1560 150
rect 2010 120 2040 150
rect 1155 60 1185 90
rect 1260 60 1290 90
rect 1800 60 1830 90
rect 1905 60 1935 90
<< metal1 >>
rect 120 1080 180 1140
rect 240 1080 300 1140
rect 360 1080 420 1140
rect 480 1080 540 1140
rect 600 1080 660 1140
rect 720 1080 780 1140
rect 840 1080 900 1140
rect 960 1080 1020 1140
rect 1080 1080 1140 1140
rect 1200 1080 1260 1140
rect 1320 1080 1380 1140
rect 1440 1080 1500 1140
rect 120 60 180 120
<< labels >>
rlabel pdiff 1562 347 1562 347 3 #22
rlabel pdiff 1427 347 1427 347 3 Vdd
rlabel pdiff 1292 347 1292 347 3 #9
rlabel poly 1502 317 1502 317 3 out
rlabel poly 1397 317 1397 317 3 in(0)
rlabel poly 1262 317 1262 317 3 in(2)
rlabel ndiff 1562 152 1562 152 3 #22
rlabel poly 1502 242 1502 242 3 out
rlabel poly 1157 317 1157 317 3 in(6)
rlabel pdiff 647 347 647 347 3 out
rlabel ndiff 1427 152 1427 152 3 GND
rlabel poly 1397 242 1397 242 3 in(0)
rlabel poly 722 317 722 317 3 in(7)
rlabel poly 617 317 617 317 3 in(5)
rlabel ndiff 1292 92 1292 92 3 out
rlabel poly 1262 242 1262 242 3 in(2)
rlabel poly 542 317 542 317 3 in(4)
rlabel poly 1157 242 1157 242 3 in(8)
rlabel poly 467 317 467 317 3 in(2)
rlabel ndiff 1052 152 1052 152 3 GND
rlabel poly 722 242 722 242 3 Vdd
rlabel poly 332 317 332 317 3 in(3)
rlabel ndiff 647 152 647 152 3 #24
rlabel pdiff 227 347 227 347 3 #9
rlabel poly 197 317 197 317 3 in(1)
rlabel pdiff 122 347 122 347 3 #10
rlabel pdiff 2297 347 2297 347 3 Vdd
rlabel poly 2087 317 2087 317 3 GND
rlabel ndiff 2042 152 2042 152 3 #24
rlabel poly 2012 242 2012 242 3 #22
rlabel poly 2012 317 2012 317 3 #22
rlabel ndiff 1937 92 1937 92 3 out
rlabel pdiff 1937 347 1937 347 3 out
rlabel poly 1907 242 1907 242 3 in(2)
rlabel poly 1907 317 1907 317 3 in(2)
rlabel pdiff 1832 347 1832 347 3 #10
rlabel poly 1802 242 1802 242 3 in(9)
rlabel ndiff 1727 92 1727 92 3 GND
rlabel metal1 1442 1082 1442 1082 3 GND
port 1 e
rlabel metal1 1322 1082 1322 1082 3 Vdd
port 2 e
rlabel metal1 1202 1082 1202 1082 3 in(9)
port 3 e
rlabel metal1 1082 1082 1082 1082 3 in(8)
port 4 e
rlabel metal1 962 1082 962 1082 3 in(7)
port 5 e
rlabel metal1 842 1082 842 1082 3 in(6)
port 6 e
rlabel metal1 722 1082 722 1082 3 in(5)
port 7 e
rlabel metal1 602 1082 602 1082 3 in(4)
port 8 e
rlabel metal1 482 1082 482 1082 3 in(3)
port 9 e
rlabel metal1 362 1082 362 1082 3 in(2)
port 10 e
rlabel metal1 242 1082 242 1082 3 in(1)
port 11 e
rlabel metal1 122 62 122 62 3 out
port 12 e
rlabel metal1 122 1082 122 1082 3 in(0)
port 13 e
<< end >>
