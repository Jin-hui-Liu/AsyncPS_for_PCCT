magic
tech sky130A
timestamp 1753015925
<< checkpaint >>
rect 57870 530370 509130 556380
rect 57870 458370 509130 511380
rect 57870 361620 509130 428130
rect 57870 255870 509130 322380
rect 57870 168120 509130 227880
rect 57870 62370 509130 128880
<< nwell >>
rect 58500 531000 508500 555750
rect 58500 459000 508500 510750
rect 58500 362250 508500 427500
rect 58500 256500 508500 321750
rect 58500 168750 508500 227250
rect 58500 63000 508500 128250
<< labels >>
rlabel nwell 58501 63001 58501 63001 3 Vdd
rlabel nwell 58501 168751 58501 168751 3 Vdd
rlabel nwell 58501 256501 58501 256501 3 Vdd
rlabel nwell 58501 362251 58501 362251 3 Vdd
rlabel nwell 58501 459001 58501 459001 3 Vdd
rlabel nwell 58501 531001 58501 531001 3 Vdd
<< end >>
