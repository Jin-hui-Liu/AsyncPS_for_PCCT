magic
tech sky130A
magscale 1 2
timestamp 1753296582
<< nwell >>
rect 180 615 945 975
rect 180 435 1320 615
rect 1575 435 1845 975
<< nmos >>
rect 195 60 225 360
rect 300 60 330 360
rect 405 270 435 360
rect 510 270 570 360
rect 915 270 945 360
rect 990 270 1320 360
rect 1425 60 1455 360
rect 1695 60 1725 360
<< pmos >>
rect 300 480 330 930
rect 405 480 435 930
rect 510 480 570 630
rect 810 480 840 930
rect 915 480 945 570
rect 990 480 1200 570
rect 1695 480 1725 930
<< ndiff >>
rect 120 330 195 360
rect 120 285 135 330
rect 180 285 195 330
rect 120 60 195 285
rect 225 60 300 360
rect 330 330 405 360
rect 330 285 345 330
rect 390 285 405 330
rect 330 270 405 285
rect 435 330 510 360
rect 435 285 450 330
rect 495 285 510 330
rect 435 270 510 285
rect 570 345 645 360
rect 570 300 585 345
rect 630 300 645 345
rect 570 270 645 300
rect 840 345 915 360
rect 840 300 855 345
rect 900 300 915 345
rect 840 270 915 300
rect 945 270 990 360
rect 1320 330 1425 360
rect 1320 285 1350 330
rect 1395 285 1425 330
rect 1320 270 1425 285
rect 330 60 390 270
rect 450 180 495 270
rect 855 105 900 270
rect 1365 60 1425 270
rect 1455 150 1530 360
rect 1455 105 1470 150
rect 1515 105 1530 150
rect 1455 60 1530 105
rect 1620 330 1695 360
rect 1620 285 1635 330
rect 1680 285 1695 330
rect 1620 60 1695 285
rect 1725 150 1800 360
rect 1725 105 1740 150
rect 1785 105 1800 150
rect 1725 60 1800 105
<< pdiff >>
rect 225 900 300 930
rect 225 855 240 900
rect 285 855 300 900
rect 225 480 300 855
rect 330 480 405 930
rect 435 630 495 930
rect 735 825 810 930
rect 735 780 750 825
rect 795 780 810 825
rect 435 555 510 630
rect 435 510 450 555
rect 495 510 510 555
rect 435 480 510 510
rect 570 540 645 630
rect 570 495 585 540
rect 630 495 645 540
rect 570 480 645 495
rect 735 480 810 780
rect 840 570 900 930
rect 1620 900 1695 930
rect 1620 855 1635 900
rect 1680 855 1695 900
rect 840 540 915 570
rect 840 495 855 540
rect 900 495 915 540
rect 840 480 915 495
rect 945 480 990 570
rect 1200 540 1275 570
rect 1200 495 1215 540
rect 1260 495 1275 540
rect 1200 480 1275 495
rect 1620 480 1695 855
rect 1725 825 1800 930
rect 1725 780 1740 825
rect 1785 780 1800 825
rect 1725 480 1800 780
<< ndiffc >>
rect 135 285 180 330
rect 345 285 390 330
rect 450 285 495 330
rect 585 300 630 345
rect 855 300 900 345
rect 1350 285 1395 330
rect 1470 105 1515 150
rect 1635 285 1680 330
rect 1740 105 1785 150
<< pdiffc >>
rect 240 855 285 900
rect 750 780 795 825
rect 450 510 495 555
rect 585 495 630 540
rect 1635 855 1680 900
rect 855 495 900 540
rect 1215 495 1260 540
rect 1740 780 1785 825
<< poly >>
rect 195 1050 330 1080
rect 195 1005 225 1050
rect 270 1005 330 1050
rect 195 975 330 1005
rect 300 930 330 975
rect 405 1050 540 1080
rect 405 1005 465 1050
rect 510 1005 540 1050
rect 405 975 540 1005
rect 780 1035 885 1065
rect 780 990 810 1035
rect 855 990 885 1035
rect 405 930 435 975
rect 780 960 885 990
rect 1650 1050 1755 1080
rect 1650 1005 1680 1050
rect 1725 1005 1755 1050
rect 1650 975 1755 1005
rect 810 930 840 960
rect 1695 930 1725 975
rect 510 630 570 660
rect 930 720 1035 750
rect 930 675 960 720
rect 1005 675 1035 720
rect 915 645 1035 675
rect 1080 675 1185 705
rect 915 570 945 645
rect 1080 630 1110 675
rect 1155 630 1185 675
rect 1080 600 1185 630
rect 990 570 1200 600
rect 300 450 330 480
rect 195 360 225 390
rect 300 360 330 390
rect 405 360 435 480
rect 510 360 570 480
rect 810 450 840 480
rect 915 360 945 480
rect 990 450 1200 480
rect 990 360 1320 390
rect 1425 360 1455 390
rect 1695 360 1725 480
rect 405 240 435 270
rect 510 195 570 270
rect 510 165 645 195
rect 510 120 570 165
rect 615 120 645 165
rect 510 90 645 120
rect 915 240 945 270
rect 990 240 1320 270
rect 1200 210 1305 240
rect 1200 165 1230 210
rect 1275 165 1305 210
rect 1200 135 1305 165
rect 195 30 225 60
rect 120 0 225 30
rect 120 -45 150 0
rect 195 -45 225 0
rect 120 -75 225 -45
rect 300 30 330 60
rect 1425 30 1455 60
rect 1695 30 1725 60
rect 300 0 405 30
rect 300 -45 330 0
rect 375 -45 405 0
rect 300 -75 405 -45
rect 1380 0 1485 30
rect 1380 -45 1410 0
rect 1455 -45 1485 0
rect 1380 -75 1485 -45
<< polycont >>
rect 225 1005 270 1050
rect 465 1005 510 1050
rect 810 990 855 1035
rect 1680 1005 1725 1050
rect 960 675 1005 720
rect 1110 630 1155 675
rect 570 120 615 165
rect 1230 165 1275 210
rect 150 -45 195 0
rect 330 -45 375 0
rect 1410 -45 1455 0
<< locali >>
rect 195 1050 300 1080
rect 195 1005 225 1050
rect 270 1005 300 1050
rect 195 975 300 1005
rect 435 1050 540 1080
rect 435 1005 465 1050
rect 510 1005 540 1050
rect 435 975 540 1005
rect 780 1035 885 1065
rect 780 990 810 1035
rect 855 990 885 1035
rect 780 960 885 990
rect 1650 1050 1755 1080
rect 1650 1005 1680 1050
rect 1725 1005 1755 1050
rect 1650 975 1755 1005
rect 240 900 285 930
rect 1635 900 1680 930
rect 240 825 285 855
rect 750 825 795 855
rect 1635 825 1680 855
rect 1740 825 1785 855
rect 750 750 795 780
rect 1740 750 1785 780
rect 930 720 1035 750
rect 930 675 960 720
rect 1005 675 1035 720
rect 930 645 1035 675
rect 1080 675 1185 705
rect 450 555 495 585
rect 450 480 495 510
rect 585 540 630 630
rect 1080 630 1110 675
rect 1155 630 1185 675
rect 1080 600 1185 630
rect 135 330 180 360
rect 135 255 180 285
rect 345 330 390 360
rect 345 150 390 285
rect 450 330 495 360
rect 450 225 495 285
rect 585 345 630 495
rect 585 270 630 300
rect 855 540 900 570
rect 855 345 900 495
rect 540 165 645 195
rect 540 120 570 165
rect 615 120 645 165
rect 540 90 645 120
rect 855 150 900 300
rect 1080 225 1125 600
rect 1215 540 1260 570
rect 1215 240 1260 495
rect 1350 330 1395 360
rect 1200 210 1305 240
rect 1200 165 1230 210
rect 1275 165 1305 210
rect 1350 225 1395 285
rect 1635 330 1680 360
rect 1635 255 1680 285
rect 1350 165 1395 180
rect 1200 135 1305 165
rect 1470 150 1515 180
rect 1470 75 1515 105
rect 1740 150 1785 180
rect 1740 75 1785 105
rect 120 0 225 30
rect 120 -45 150 0
rect 195 -45 225 0
rect 120 -75 225 -45
rect 300 0 405 30
rect 300 -45 330 0
rect 375 -45 405 0
rect 300 -75 405 -45
rect 1380 0 1485 30
rect 1380 -45 1410 0
rect 1455 -45 1485 0
rect 1380 -75 1485 -45
<< viali >>
rect 225 1005 270 1050
rect 465 1005 510 1050
rect 810 990 855 1035
rect 1680 1005 1725 1050
rect 240 855 285 900
rect 1635 855 1680 900
rect 750 780 795 825
rect 1740 780 1785 825
rect 960 675 1005 720
rect 585 630 630 675
rect 135 285 180 330
rect 450 180 495 225
rect 345 105 390 150
rect 570 120 615 165
rect 1215 495 1260 540
rect 1080 180 1125 225
rect 855 105 900 150
rect 1635 285 1680 330
rect 1350 180 1395 225
rect 1470 105 1515 150
rect 1740 105 1785 150
rect 150 -45 195 0
rect 330 -45 375 0
rect 1410 -45 1455 0
<< metal1 >>
rect 210 1050 285 1065
rect 210 1005 225 1050
rect 270 1005 285 1050
rect 210 990 285 1005
rect 450 1050 525 1065
rect 1665 1050 1740 1065
rect 450 1005 465 1050
rect 510 1005 525 1050
rect 450 990 525 1005
rect 795 1035 870 1050
rect 795 990 810 1035
rect 855 990 870 1035
rect 1665 1005 1680 1050
rect 1725 1005 1740 1050
rect 1665 990 1740 1005
rect 795 975 870 990
rect 225 900 1695 915
rect 225 855 240 900
rect 285 885 1635 900
rect 285 855 300 885
rect 225 840 300 855
rect 1620 855 1635 885
rect 1680 855 1695 900
rect 1620 840 1695 855
rect 735 825 810 840
rect 735 780 750 825
rect 795 810 810 825
rect 1725 825 1800 840
rect 1725 810 1740 825
rect 795 780 1740 810
rect 1785 780 1800 825
rect 735 765 810 780
rect 1725 765 1800 780
rect 945 720 1020 735
rect 945 690 960 720
rect 570 675 960 690
rect 1005 675 1020 720
rect 570 630 585 675
rect 630 660 1020 675
rect 630 630 645 660
rect 570 615 645 630
rect 435 540 510 570
rect 1200 540 1275 555
rect 435 510 1215 540
rect 435 495 510 510
rect 1200 495 1215 510
rect 1260 495 1275 540
rect 1200 480 1275 495
rect 120 330 1695 345
rect 120 285 135 330
rect 180 315 1635 330
rect 180 285 195 315
rect 120 270 195 285
rect 1620 285 1635 315
rect 1680 285 1695 330
rect 1620 270 1695 285
rect 435 225 1410 240
rect 435 180 450 225
rect 495 210 1080 225
rect 495 180 510 210
rect 1065 180 1080 210
rect 1125 210 1350 225
rect 1125 180 1140 210
rect 435 165 510 180
rect 555 165 630 180
rect 1065 165 1140 180
rect 1335 180 1350 210
rect 1395 180 1410 225
rect 1335 165 1410 180
rect 330 150 405 165
rect 330 105 345 150
rect 390 135 405 150
rect 555 135 570 165
rect 390 120 570 135
rect 615 135 630 165
rect 840 150 915 165
rect 840 135 855 150
rect 615 120 855 135
rect 390 105 855 120
rect 900 105 915 150
rect 330 90 405 105
rect 840 90 915 105
rect 1455 150 1800 165
rect 1455 105 1470 150
rect 1515 135 1740 150
rect 1515 105 1530 135
rect 1455 90 1530 105
rect 1725 105 1740 135
rect 1785 105 1800 150
rect 1725 90 1800 105
rect 135 0 210 15
rect 135 -45 150 0
rect 195 -45 210 0
rect 135 -60 210 -45
rect 315 0 390 15
rect 315 -45 330 0
rect 375 -45 390 0
rect 315 -60 390 -45
rect 1395 0 1470 15
rect 1395 -45 1410 0
rect 1455 -45 1470 0
rect 1395 -60 1470 -45
<< labels >>
flabel ndiff 360 60 360 60 1 FreeSerif 120 0 0 0 out
flabel ndiff 1485 60 1485 60 1 FreeSerif 120 0 0 0 #6
flabel ndiff 1650 60 1650 60 1 FreeSerif 120 0 0 0 #5
flabel ndiff 1755 60 1755 60 1 FreeSerif 120 0 0 0 #6
flabel ndiff 465 270 465 270 1 FreeSerif 120 0 0 0 GND
flabel ndiff 600 270 600 270 1 FreeSerif 120 0 0 0 #16
flabel poly 510 405 510 405 3 FreeSerif 120 0 0 0 out
flabel poly 405 405 405 405 3 FreeSerif 120 0 0 0 in(0)
flabel poly 195 375 195 375 3 FreeSerif 120 0 0 0 in(5)
flabel poly 300 375 300 375 3 FreeSerif 120 0 0 0 in(6)
flabel ndiff 870 270 870 270 1 FreeSerif 120 0 0 0 out
flabel poly 1020 375 1020 375 3 FreeSerif 120 0 0 0 Vdd
flabel poly 915 405 915 405 3 FreeSerif 120 0 0 0 #16
flabel poly 810 465 810 465 3 FreeSerif 120 0 0 0 in(3)
flabel poly 1020 465 1020 465 3 FreeSerif 120 0 0 0 GND
flabel ndiff 1335 315 1335 315 3 FreeSerif 120 0 0 0 GND
flabel poly 1695 420 1695 420 3 FreeSerif 120 0 0 0 in(2)
flabel poly 1425 375 1425 375 3 FreeSerif 120 0 0 0 in(4)
flabel pdiff 1770 480 1770 480 1 FreeSerif 120 0 0 0 #11
flabel pdiff 1665 480 1665 480 1 FreeSerif 120 0 0 0 #12
flabel pdiff 1230 495 1230 495 3 FreeSerif 120 0 0 0 Vdd
flabel pdiff 855 495 855 495 1 FreeSerif 120 0 0 0 out
flabel pdiff 750 495 750 495 1 FreeSerif 120 0 0 0 #11
flabel pdiff 600 480 600 480 1 FreeSerif 120 0 0 0 #16
flabel pdiff 465 480 465 480 1 FreeSerif 120 0 0 0 Vdd
flabel poly 300 465 300 465 3 FreeSerif 120 0 0 0 in(1)
flabel pdiff 255 480 255 480 1 FreeSerif 120 0 0 0 #12
flabel ndiff 150 60 150 60 1 FreeSerif 120 0 0 0 #5
flabel metal1 1095 165 1095 165 5 FreeSerif 120 0 0 0 GND
port 1 s
flabel metal1 1275 510 1275 510 3 FreeSerif 120 0 0 0 Vdd
port 2 e
flabel metal1 165 -60 165 -60 5 FreeSerif 120 0 0 0 in(5)
port 4 s
flabel metal1 345 -60 345 -60 5 FreeSerif 120 0 0 0 in(6)
port 3 s
flabel metal1 1425 -60 1425 -60 5 FreeSerif 120 0 0 0 in(4)
port 5 s
flabel metal1 1695 1065 1695 1065 1 FreeSerif 120 0 0 0 in(2)
port 7 n
flabel metal1 825 1050 825 1050 1 FreeSerif 120 0 0 0 in(3)
port 6 n
flabel metal1 495 1065 495 1065 1 FreeSerif 120 0 0 0 in(0)
port 10 n
flabel metal1 240 1065 240 1065 1 FreeSerif 120 0 0 0 in(1)
port 8 n
flabel metal1 600 105 600 105 5 FreeSerif 120 0 0 0 out
port 9 s
<< end >>
