magic
tech sky130A
magscale 1 2
timestamp 1753369762
<< nwell >>
rect 315 795 675 1095
rect 1320 795 1680 1095
rect 315 735 1680 795
rect 315 555 2085 735
<< nmos >>
rect 195 285 225 480
rect 330 75 360 480
rect 435 75 465 480
rect 540 375 570 480
rect 675 180 705 480
rect 810 390 870 480
rect 1530 330 1560 480
rect 1665 180 1695 480
rect 1935 390 1965 480
rect 2010 390 2340 480
<< pmos >>
rect 435 600 465 1050
rect 540 600 570 1050
rect 675 600 705 720
rect 810 600 870 750
rect 1110 600 1320 690
rect 1425 600 1455 1050
rect 1530 600 1560 1050
rect 1935 600 1965 690
<< ndiff >>
rect 120 450 195 480
rect 120 405 135 450
rect 180 405 195 450
rect 120 285 195 405
rect 225 285 330 480
rect 270 75 330 285
rect 360 75 435 480
rect 465 465 540 480
rect 465 420 480 465
rect 525 420 540 465
rect 465 375 540 420
rect 570 450 675 480
rect 570 405 600 450
rect 645 405 675 450
rect 570 375 675 405
rect 465 75 525 375
rect 615 180 675 375
rect 705 465 810 480
rect 705 420 735 465
rect 780 420 810 465
rect 705 390 810 420
rect 870 465 945 480
rect 870 420 885 465
rect 930 420 945 465
rect 870 390 945 420
rect 1455 450 1530 480
rect 1455 405 1470 450
rect 1515 405 1530 450
rect 705 180 765 390
rect 1455 330 1530 405
rect 1560 330 1665 480
rect 1605 180 1665 330
rect 1695 465 1770 480
rect 1695 420 1710 465
rect 1755 420 1770 465
rect 1695 180 1770 420
rect 1860 465 1935 480
rect 1860 420 1875 465
rect 1920 420 1935 465
rect 1860 390 1935 420
rect 1965 390 2010 480
rect 2340 465 2415 480
rect 2340 420 2355 465
rect 2400 420 2415 465
rect 2340 390 2415 420
<< pdiff >>
rect 360 1020 435 1050
rect 360 975 375 1020
rect 420 975 435 1020
rect 360 600 435 975
rect 465 600 540 1050
rect 570 720 630 1050
rect 750 720 810 750
rect 570 705 675 720
rect 570 660 585 705
rect 630 660 675 705
rect 570 600 675 660
rect 705 675 810 720
rect 705 630 735 675
rect 780 630 810 675
rect 705 600 810 630
rect 870 660 945 750
rect 1365 690 1425 1050
rect 870 615 885 660
rect 930 615 945 660
rect 870 600 945 615
rect 1035 675 1110 690
rect 1035 630 1050 675
rect 1095 630 1110 675
rect 1035 600 1110 630
rect 1320 675 1425 690
rect 1320 630 1350 675
rect 1395 630 1425 675
rect 1320 600 1425 630
rect 1455 600 1530 1050
rect 1560 1020 1635 1050
rect 1560 975 1575 1020
rect 1620 975 1635 1020
rect 1560 600 1635 975
rect 1860 675 1935 690
rect 1860 630 1875 675
rect 1920 630 1935 675
rect 1860 600 1935 630
rect 1965 675 2040 690
rect 1965 630 1980 675
rect 2025 630 2040 675
rect 1965 600 2040 630
<< ndiffc >>
rect 135 405 180 450
rect 480 420 525 465
rect 600 405 645 450
rect 735 420 780 465
rect 885 420 930 465
rect 1470 405 1515 450
rect 1710 420 1755 465
rect 1875 420 1920 465
rect 2355 420 2400 465
<< pdiffc >>
rect 375 975 420 1020
rect 585 660 630 705
rect 735 630 780 675
rect 885 615 930 660
rect 1050 630 1095 675
rect 1350 630 1395 675
rect 1575 975 1620 1020
rect 1875 630 1920 675
rect 1980 630 2025 675
<< poly >>
rect 360 1170 465 1200
rect 360 1125 390 1170
rect 435 1125 465 1170
rect 360 1095 465 1125
rect 435 1050 465 1095
rect 540 1170 645 1200
rect 540 1125 570 1170
rect 615 1125 645 1170
rect 540 1095 645 1125
rect 1350 1155 1455 1185
rect 1350 1110 1380 1155
rect 1425 1110 1455 1155
rect 540 1050 570 1095
rect 1350 1080 1455 1110
rect 1425 1050 1455 1080
rect 1530 1050 1560 1080
rect 810 855 915 885
rect 810 810 840 855
rect 885 810 915 855
rect 810 780 915 810
rect 810 750 870 780
rect 675 720 705 750
rect 1110 690 1320 720
rect 1935 690 1965 720
rect 2145 645 2250 675
rect 2145 600 2175 645
rect 2220 600 2250 645
rect 435 570 465 600
rect 195 480 225 510
rect 330 480 360 510
rect 435 480 465 510
rect 540 480 570 600
rect 675 480 705 600
rect 810 480 870 600
rect 1110 570 1320 600
rect 1425 570 1455 600
rect 1170 540 1275 570
rect 1170 495 1200 540
rect 1245 495 1275 540
rect 195 255 225 285
rect 120 225 225 255
rect 120 180 150 225
rect 195 180 225 225
rect 120 150 225 180
rect 540 345 570 375
rect 1170 465 1275 495
rect 1530 480 1560 600
rect 1665 480 1695 510
rect 1935 480 1965 600
rect 2145 570 2250 600
rect 2175 510 2205 570
rect 2010 480 2340 510
rect 810 360 870 390
rect 1530 255 1560 330
rect 1455 225 1560 255
rect 1455 180 1485 225
rect 1530 180 1560 225
rect 1935 345 1965 390
rect 2010 360 2340 390
rect 1860 315 1965 345
rect 1860 270 1890 315
rect 1935 270 1965 315
rect 1860 240 1965 270
rect 675 150 705 180
rect 1455 150 1560 180
rect 1665 150 1695 180
rect 675 120 780 150
rect 675 75 705 120
rect 750 75 780 120
rect 330 45 360 75
rect 255 15 360 45
rect 255 -30 285 15
rect 330 -30 360 15
rect 255 -60 360 -30
rect 435 45 465 75
rect 675 45 780 75
rect 1665 120 1770 150
rect 1665 75 1695 120
rect 1740 75 1770 120
rect 1665 45 1770 75
rect 435 15 540 45
rect 435 -30 465 15
rect 510 -30 540 15
rect 435 -60 540 -30
<< polycont >>
rect 390 1125 435 1170
rect 570 1125 615 1170
rect 1380 1110 1425 1155
rect 840 810 885 855
rect 2175 600 2220 645
rect 1200 495 1245 540
rect 150 180 195 225
rect 1485 180 1530 225
rect 1890 270 1935 315
rect 705 75 750 120
rect 285 -30 330 15
rect 1695 75 1740 120
rect 465 -30 510 15
<< locali >>
rect 360 1170 465 1200
rect 360 1125 390 1170
rect 435 1125 465 1170
rect 360 1095 465 1125
rect 540 1170 645 1200
rect 540 1125 570 1170
rect 615 1125 645 1170
rect 540 1095 645 1125
rect 1350 1155 1455 1185
rect 1350 1110 1380 1155
rect 1425 1110 1455 1155
rect 1350 1080 1455 1110
rect 375 1020 420 1050
rect 375 945 420 975
rect 1575 1020 1620 1050
rect 1575 945 1620 975
rect 810 855 915 885
rect 810 810 840 855
rect 885 810 915 855
rect 135 450 180 480
rect 135 375 180 405
rect 480 465 525 765
rect 810 780 915 810
rect 585 705 630 750
rect 585 630 630 660
rect 735 675 780 705
rect 735 600 780 630
rect 885 660 930 690
rect 480 390 525 420
rect 600 450 645 480
rect 600 375 645 405
rect 735 465 780 510
rect 735 390 780 420
rect 885 465 930 615
rect 1050 675 1095 735
rect 1050 600 1095 630
rect 1350 675 1395 705
rect 1350 600 1395 630
rect 1170 540 1275 570
rect 1170 495 1200 540
rect 1245 495 1275 540
rect 1170 465 1275 495
rect 885 330 930 420
rect 1470 450 1515 480
rect 1470 375 1515 405
rect 1710 465 1755 825
rect 1875 675 1920 735
rect 1875 600 1920 630
rect 1980 675 2025 810
rect 1980 600 2025 630
rect 2145 645 2250 675
rect 2145 600 2175 645
rect 2220 600 2250 645
rect 2145 570 2250 600
rect 1875 465 1920 495
rect 1755 420 1875 465
rect 1710 390 1755 420
rect 1875 390 1920 420
rect 2355 465 2400 540
rect 2355 390 2400 420
rect 1860 315 1965 345
rect 1860 270 1890 315
rect 1935 270 1965 315
rect 120 225 225 255
rect 120 180 150 225
rect 195 180 225 225
rect 120 150 225 180
rect 1455 225 1560 255
rect 1860 240 1965 270
rect 1455 180 1485 225
rect 1530 180 1560 225
rect 1455 150 1560 180
rect 675 120 780 150
rect 675 75 705 120
rect 750 75 780 120
rect 675 45 780 75
rect 1665 120 1770 150
rect 1665 75 1695 120
rect 1740 75 1770 120
rect 1665 45 1770 75
rect 255 15 360 45
rect 255 -30 285 15
rect 330 -30 360 15
rect 255 -60 360 -30
rect 435 15 540 45
rect 435 -30 465 15
rect 510 -30 540 15
rect 435 -60 540 -30
<< viali >>
rect 390 1125 435 1170
rect 570 1125 615 1170
rect 1380 1110 1425 1155
rect 375 975 420 1020
rect 1575 975 1620 1020
rect 840 810 885 855
rect 480 765 525 810
rect 135 405 180 450
rect 585 750 630 795
rect 1710 825 1755 870
rect 1050 735 1095 780
rect 735 630 780 675
rect 735 510 780 555
rect 600 405 645 450
rect 1350 630 1395 675
rect 1200 495 1245 540
rect 1470 405 1515 450
rect 1980 810 2025 855
rect 1875 735 1920 780
rect 2175 600 2220 645
rect 2355 540 2400 585
rect 885 285 930 330
rect 1890 270 1935 315
rect 150 180 195 225
rect 1485 180 1530 225
rect 705 75 750 120
rect 1695 75 1740 120
rect 285 -30 330 15
rect 465 -30 510 15
<< metal1 >>
rect 375 1170 450 1185
rect 375 1125 390 1170
rect 435 1125 450 1170
rect 375 1110 450 1125
rect 555 1170 630 1185
rect 555 1125 570 1170
rect 615 1125 630 1170
rect 555 1110 630 1125
rect 1365 1155 1440 1170
rect 1365 1110 1380 1155
rect 1425 1110 1440 1155
rect 1365 1095 1440 1110
rect 360 1020 1635 1035
rect 360 975 375 1020
rect 420 1005 1575 1020
rect 420 975 435 1005
rect 360 960 435 975
rect 1560 975 1575 1005
rect 1620 975 1635 1020
rect 1560 960 1635 975
rect 1695 870 1770 885
rect 825 855 1710 870
rect 825 825 840 855
rect 465 810 840 825
rect 885 840 1710 855
rect 885 810 900 840
rect 1695 825 1710 840
rect 1755 855 2040 870
rect 1755 840 1980 855
rect 1755 825 1770 840
rect 1695 810 1770 825
rect 1965 810 1980 840
rect 2025 810 2040 855
rect 465 765 480 810
rect 525 795 900 810
rect 1965 795 2040 810
rect 525 765 540 795
rect 465 750 540 765
rect 570 750 585 795
rect 630 750 645 795
rect 570 735 645 750
rect 1035 780 1110 795
rect 1860 780 1935 795
rect 1035 735 1050 780
rect 1095 750 1875 780
rect 1095 735 1110 750
rect 1035 720 1110 735
rect 1860 735 1875 750
rect 1920 735 1935 780
rect 1860 720 1935 735
rect 720 675 795 690
rect 720 630 735 675
rect 780 645 795 675
rect 1335 675 1410 690
rect 1335 645 1350 675
rect 780 630 1350 645
rect 1395 645 1410 675
rect 2160 645 2235 660
rect 1395 630 2175 645
rect 720 615 2175 630
rect 2160 600 2175 615
rect 2220 600 2235 645
rect 2160 585 2235 600
rect 2340 585 2415 600
rect 720 555 795 570
rect 2340 555 2355 585
rect 720 510 735 555
rect 780 540 2355 555
rect 2400 540 2415 585
rect 780 525 1200 540
rect 780 510 795 525
rect 720 495 795 510
rect 1185 495 1200 525
rect 1245 525 2415 540
rect 1245 495 1260 525
rect 1185 480 1260 495
rect 120 450 195 465
rect 120 405 135 450
rect 180 420 195 450
rect 585 450 660 465
rect 585 420 600 450
rect 180 405 600 420
rect 645 420 660 450
rect 1455 450 1530 465
rect 1455 420 1470 450
rect 645 405 1470 420
rect 1515 405 1530 450
rect 120 390 1530 405
rect 870 330 945 345
rect 870 285 885 330
rect 930 315 1950 330
rect 930 300 1890 315
rect 930 285 945 300
rect 870 270 945 285
rect 1875 270 1890 300
rect 1935 270 1950 315
rect 1875 255 1950 270
rect 135 225 1545 240
rect 135 180 150 225
rect 195 210 1485 225
rect 195 180 210 210
rect 135 165 210 180
rect 1470 180 1485 210
rect 1530 180 1545 225
rect 1470 165 1545 180
rect 690 120 765 135
rect 690 75 705 120
rect 750 75 765 120
rect 690 60 765 75
rect 1680 120 1755 135
rect 1680 75 1695 120
rect 1740 75 1755 120
rect 1680 60 1755 75
rect 270 15 345 30
rect 270 -30 285 15
rect 330 -30 345 15
rect 270 -45 345 -30
rect 450 15 525 30
rect 450 -30 465 15
rect 510 -30 525 15
rect 450 -45 525 -30
<< labels >>
flabel poly 195 495 195 495 3 FreeSerif 120 0 0 0 in(2)
flabel poly 330 495 330 495 3 FreeSerif 120 0 0 0 in(6)
flabel poly 435 495 435 495 3 FreeSerif 120 0 0 0 in(7)
flabel poly 435 585 435 585 3 FreeSerif 120 0 0 0 in(3)
flabel poly 540 540 540 540 3 FreeSerif 120 0 0 0 in(4)
flabel poly 675 540 675 540 3 FreeSerif 120 0 0 0 in(0)
flabel poly 810 540 810 540 3 FreeSerif 120 0 0 0 out
flabel poly 1140 585 1140 585 3 FreeSerif 120 0 0 0 GND
flabel poly 1425 585 1425 585 3 FreeSerif 120 0 0 0 in(1)
flabel poly 1530 540 1530 540 3 FreeSerif 120 0 0 0 in(2)
flabel poly 1665 495 1665 495 3 FreeSerif 120 0 0 0 in(5)
flabel poly 1935 540 1935 540 3 FreeSerif 120 0 0 0 #18
flabel poly 2040 495 2040 495 3 FreeSerif 120 0 0 0 Vdd
flabel pdiff 405 600 405 600 1 FreeSerif 120 0 0 0 #14
flabel pdiff 630 600 630 600 1 FreeSerif 120 0 0 0 out
flabel pdiff 765 600 765 600 1 FreeSerif 120 0 0 0 Vdd
flabel pdiff 915 600 915 600 1 FreeSerif 120 0 0 0 #18
flabel pdiff 1080 600 1080 600 1 FreeSerif 120 0 0 0 #19
flabel pdiff 1380 600 1380 600 1 FreeSerif 120 0 0 0 Vdd
flabel pdiff 1605 600 1605 600 1 FreeSerif 120 0 0 0 #14
flabel pdiff 1905 600 1905 600 1 FreeSerif 120 0 0 0 #19
flabel pdiff 2010 600 2010 600 1 FreeSerif 120 0 0 0 out
flabel ndiff 1905 390 1905 390 1 FreeSerif 120 0 0 0 out
flabel ndiff 2385 390 2385 390 1 FreeSerif 120 0 0 0 GND
flabel ndiff 1500 330 1500 330 1 FreeSerif 120 0 0 0 #3
flabel ndiff 1740 180 1740 180 1 FreeSerif 120 0 0 0 out
flabel ndiff 915 390 915 390 1 FreeSerif 120 0 0 0 #18
flabel ndiff 720 195 720 195 3 FreeSerif 120 0 0 0 GND
flabel ndiff 615 375 615 375 1 FreeSerif 120 0 0 0 #3
flabel ndiff 495 75 495 75 1 FreeSerif 120 0 0 0 out
flabel ndiff 150 285 150 285 1 FreeSerif 120 0 0 0 #3
flabel metal1 1215 480 1215 480 5 FreeSerif 120 0 0 0 GND
port 1 s
flabel metal1 2190 660 2190 660 1 FreeSerif 120 0 0 0 Vdd
port 2 n
flabel metal1 495 -45 495 -45 5 FreeSerif 120 0 0 0 in(7)
port 3 s
flabel metal1 300 -45 300 -45 5 FreeSerif 120 0 0 0 in(6)
port 4 s
flabel metal1 1725 60 1725 60 5 FreeSerif 120 0 0 0 in(5)
port 5 s
flabel metal1 600 1185 600 1185 1 FreeSerif 120 0 0 0 in(4)
port 6 n
flabel metal1 405 1185 405 1185 1 FreeSerif 120 0 0 0 in(3)
port 7 n
flabel metal1 1485 165 1485 165 5 FreeSerif 120 0 0 0 in(2)
port 8 s
flabel metal1 1395 1170 1395 1170 1 FreeSerif 120 0 0 0 in(1)
port 9 n
flabel metal1 855 870 855 870 1 FreeSerif 120 0 0 0 out
port 10 n
flabel metal1 735 60 735 60 5 FreeSerif 120 0 0 0 in(0)
port 11 s
<< end >>
